library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;


package FACE_DETECTION_PCK is

constant IMG_WIDTH : integer := 128;
constant IMG_HEIGHT: integer :=64;

type STAGE_NF is array (0 to 24 ) of integer;
type FEATURE_NR  is array (0 to 2912) of integer;

constant SNF : STAGE_NF := (0 => 9,
1 => 16,
2 => 27,
3 => 32,
4 => 52,
5 => 53,
6 => 62,
7 => 72,
8 => 83,
9 => 91,
10 => 99,
11 => 115,
12 => 127,
13 => 135,
14 => 136,
15 => 137,
16 => 159,
17 => 155,
18 => 169,
19 => 196,
20 => 197,
21 => 181,
22 => 199,
23 => 211,
24 => 200); -- TODO:

constant FNR : FEATURE_NR := (
0 => 2,
1 => 2,
2 => 2,
3 => 2,
4 => 2,
5 => 2,
6 => 2,
7 => 2,
8 => 2,
9 => 2,
10 => 2,
11 => 2,
12 => 2,
13 => 2,
14 => 2,
15 => 2,
16 => 2,
17 => 2,
18 => 2,
19 => 2,
20 => 2,
21 => 2,
22 => 2,
23 => 2,
24 => 2,
25 => 2,
26 => 2,
27 => 2,
28 => 2,
29 => 2,
30 => 2,
31 => 2,
32 => 2,
33 => 2,
34 => 2,
35 => 3,
36 => 2,
37 => 2,
38 => 2,
39 => 2,
40 => 2,
41 => 2,
42 => 2,
43 => 2,
44 => 2,
45 => 2,
46 => 2,
47 => 2,
48 => 3,
49 => 2,
50 => 2,
51 => 2,
52 => 2,
53 => 2,
54 => 2,
55 => 2,
56 => 3,
57 => 2,
58 => 2,
59 => 2,
60 => 2,
61 => 2,
62 => 3,
63 => 2,
64 => 2,
65 => 2,
66 => 2,
67 => 2,
68 => 2,
69 => 2,
70 => 3,
71 => 2,
72 => 2,
73 => 2,
74 => 2,
75 => 3,
76 => 3,
77 => 2,
78 => 2,
79 => 2,
80 => 2,
81 => 2,
82 => 2,
83 => 2,
84 => 2,
85 => 2,
86 => 2,
87 => 2,
88 => 2,
89 => 2,
90 => 2,
91 => 2,
92 => 2,
93 => 2,
94 => 2,
95 => 2,
96 => 2,
97 => 2,
98 => 2,
99 => 2,
100 => 2,
101 => 2,
102 => 2,
103 => 2,
104 => 2,
105 => 3,
106 => 2,
107 => 2,
108 => 2,
109 => 3,
110 => 3,
111 => 2,
112 => 2,
113 => 2,
114 => 2,
115 => 2,
116 => 2,
117 => 2,
118 => 3,
119 => 2,
120 => 3,
121 => 3,
122 => 3,
123 => 2,
124 => 2,
125 => 2,
126 => 2,
127 => 2,
128 => 2,
129 => 2,
130 => 2,
131 => 2,
132 => 2,
133 => 2,
134 => 2,
135 => 2,
136 => 2,
137 => 2,
138 => 2,
139 => 2,
140 => 2,
141 => 2,
142 => 2,
143 => 2,
144 => 2,
145 => 2,
146 => 2,
147 => 2,
148 => 2,
149 => 2,
150 => 2,
151 => 2,
152 => 3,
153 => 2,
154 => 2,
155 => 2,
156 => 2,
157 => 2,
158 => 2,
159 => 2,
160 => 3,
161 => 2,
162 => 2,
163 => 2,
164 => 3,
165 => 2,
166 => 2,
167 => 2,
168 => 2,
169 => 2,
170 => 2,
171 => 2,
172 => 2,
173 => 2,
174 => 2,
175 => 2,
176 => 3,
177 => 3,
178 => 2,
179 => 2,
180 => 2,
181 => 2,
182 => 2,
183 => 2,
184 => 2,
185 => 2,
186 => 2,
187 => 3,
188 => 2,
189 => 2,
190 => 2,
191 => 2,
192 => 2,
193 => 2,
194 => 2,
195 => 2,
196 => 2,
197 => 2,
198 => 2,
199 => 2,
200 => 2,
201 => 2,
202 => 3,
203 => 2,
204 => 2,
205 => 2,
206 => 3,
207 => 3,
208 => 2,
209 => 2,
210 => 2,
211 => 2,
212 => 2,
213 => 2,
214 => 2,
215 => 3,
216 => 2,
217 => 3,
218 => 2,
219 => 2,
220 => 2,
221 => 2,
222 => 2,
223 => 3,
224 => 3,
225 => 2,
226 => 2,
227 => 2,
228 => 2,
229 => 2,
230 => 3,
231 => 2,
232 => 2,
233 => 2,
234 => 3,
235 => 3,
236 => 2,
237 => 2,
238 => 2,
239 => 2,
240 => 2,
241 => 3,
242 => 3,
243 => 2,
244 => 2,
245 => 2,
246 => 2,
247 => 2,
248 => 3,
249 => 3,
250 => 2,
251 => 2,
252 => 2,
253 => 2,
254 => 2,
255 => 3,
256 => 2,
257 => 2,
258 => 2,
259 => 2,
260 => 2,
261 => 3,
262 => 2,
263 => 2,
264 => 2,
265 => 2,
266 => 2,
267 => 2,
268 => 2,
269 => 2,
270 => 2,
271 => 2,
272 => 2,
273 => 2,
274 => 2,
275 => 2,
276 => 2,
277 => 2,
278 => 2,
279 => 2,
280 => 2,
281 => 2,
282 => 2,
283 => 2,
284 => 2,
285 => 2,
286 => 2,
287 => 2,
288 => 3,
289 => 2,
290 => 2,
291 => 3,
292 => 2,
293 => 2,
294 => 2,
295 => 2,
296 => 2,
297 => 2,
298 => 2,
299 => 2,
300 => 2,
301 => 2,
302 => 2,
303 => 2,
304 => 2,
305 => 2,
306 => 2,
307 => 2,
308 => 2,
309 => 2,
310 => 2,
311 => 2,
312 => 2,
313 => 2,
314 => 2,
315 => 2,
316 => 2,
317 => 3,
318 => 3,
319 => 3,
320 => 2,
321 => 2,
322 => 2,
323 => 2,
324 => 2,
325 => 2,
326 => 2,
327 => 3,
328 => 2,
329 => 2,
330 => 2,
331 => 2,
332 => 2,
333 => 2,
334 => 2,
335 => 2,
336 => 3,
337 => 3,
338 => 2,
339 => 2,
340 => 2,
341 => 2,
342 => 2,
343 => 2,
344 => 2,
345 => 2,
346 => 2,
347 => 2,
348 => 2,
349 => 2,
350 => 2,
351 => 2,
352 => 2,
353 => 2,
354 => 2,
355 => 2,
356 => 2,
357 => 2,
358 => 2,
359 => 3,
360 => 3,
361 => 3,
362 => 3,
363 => 3,
364 => 2,
365 => 2,
366 => 3,
367 => 3,
368 => 2,
369 => 2,
370 => 2,
371 => 2,
372 => 2,
373 => 3,
374 => 3,
375 => 3,
376 => 2,
377 => 2,
378 => 2,
379 => 2,
380 => 2,
381 => 2,
382 => 2,
383 => 2,
384 => 2,
385 => 2,
386 => 2,
387 => 2,
388 => 2,
389 => 2,
390 => 2,
391 => 2,
392 => 2,
393 => 2,
394 => 2,
395 => 2,
396 => 2,
397 => 2,
398 => 2,
399 => 2,
400 => 2,
401 => 2,
402 => 2,
403 => 2,
404 => 2,
405 => 2,
406 => 2,
407 => 2,
408 => 2,
409 => 2,
410 => 2,
411 => 2,
412 => 3,
413 => 2,
414 => 2,
415 => 3,
416 => 3,
417 => 2,
418 => 2,
419 => 2,
420 => 2,
421 => 2,
422 => 2,
423 => 2,
424 => 2,
425 => 2,
426 => 2,
427 => 2,
428 => 2,
429 => 2,
430 => 2,
431 => 2,
432 => 2,
433 => 2,
434 => 2,
435 => 2,
436 => 2,
437 => 2,
438 => 2,
439 => 2,
440 => 2,
441 => 2,
442 => 2,
443 => 2,
444 => 3,
445 => 2,
446 => 2,
447 => 2,
448 => 2,
449 => 2,
450 => 2,
451 => 3,
452 => 2,
453 => 3,
454 => 3,
455 => 2,
456 => 2,
457 => 2,
458 => 2,
459 => 3,
460 => 3,
461 => 3,
462 => 2,
463 => 3,
464 => 3,
465 => 2,
466 => 2,
467 => 2,
468 => 2,
469 => 2,
470 => 2,
471 => 2,
472 => 2,
473 => 3,
474 => 2,
475 => 2,
476 => 2,
477 => 2,
478 => 3,
479 => 2,
480 => 2,
481 => 3,
482 => 2,
483 => 2,
484 => 2,
485 => 2,
486 => 2,
487 => 2,
488 => 2,
489 => 2,
490 => 3,
491 => 2,
492 => 2,
493 => 2,
494 => 2,
495 => 2,
496 => 2,
497 => 2,
498 => 2,
499 => 2,
500 => 2,
501 => 2,
502 => 2,
503 => 2,
504 => 2,
505 => 2,
506 => 2,
507 => 2,
508 => 2,
509 => 2,
510 => 2,
511 => 2,
512 => 2,
513 => 2,
514 => 2,
515 => 2,
516 => 2,
517 => 2,
518 => 2,
519 => 2,
520 => 3,
521 => 3,
522 => 2,
523 => 2,
524 => 2,
525 => 3,
526 => 2,
527 => 2,
528 => 2,
529 => 3,
530 => 2,
531 => 2,
532 => 2,
533 => 2,
534 => 2,
535 => 2,
536 => 2,
537 => 2,
538 => 2,
539 => 2,
540 => 2,
541 => 2,
542 => 3,
543 => 2,
544 => 2,
545 => 2,
546 => 3,
547 => 2,
548 => 3,
549 => 3,
550 => 2,
551 => 2,
552 => 2,
553 => 2,
554 => 3,
555 => 2,
556 => 2,
557 => 2,
558 => 2,
559 => 3,
560 => 2,
561 => 2,
562 => 2,
563 => 2,
564 => 2,
565 => 2,
566 => 2,
567 => 2,
568 => 2,
569 => 2,
570 => 2,
571 => 2,
572 => 2,
573 => 2,
574 => 2,
575 => 2,
576 => 2,
577 => 2,
578 => 2,
579 => 2,
580 => 2,
581 => 2,
582 => 2,
583 => 2,
584 => 2,
585 => 2,
586 => 2,
587 => 3,
588 => 3,
589 => 2,
590 => 2,
591 => 3,
592 => 3,
593 => 2,
594 => 3,
595 => 3,
596 => 2,
597 => 2,
598 => 2,
599 => 2,
600 => 2,
601 => 2,
602 => 2,
603 => 2,
604 => 2,
605 => 2,
606 => 2,
607 => 2,
608 => 2,
609 => 2,
610 => 2,
611 => 2,
612 => 2,
613 => 2,
614 => 2,
615 => 2,
616 => 2,
617 => 2,
618 => 2,
619 => 2,
620 => 2,
621 => 2,
622 => 2,
623 => 2,
624 => 3,
625 => 3,
626 => 2,
627 => 2,
628 => 2,
629 => 2,
630 => 2,
631 => 2,
632 => 2,
633 => 2,
634 => 2,
635 => 2,
636 => 2,
637 => 2,
638 => 2,
639 => 2,
640 => 2,
641 => 2,
642 => 2,
643 => 2,
644 => 2,
645 => 2,
646 => 2,
647 => 2,
648 => 2,
649 => 2,
650 => 2,
651 => 2,
652 => 2,
653 => 2,
654 => 2,
655 => 3,
656 => 2,
657 => 2,
658 => 2,
659 => 3,
660 => 2,
661 => 2,
662 => 2,
663 => 2,
664 => 2,
665 => 3,
666 => 3,
667 => 2,
668 => 2,
669 => 2,
670 => 2,
671 => 2,
672 => 2,
673 => 2,
674 => 2,
675 => 3,
676 => 2,
677 => 2,
678 => 3,
679 => 3,
680 => 3,
681 => 2,
682 => 2,
683 => 3,
684 => 2,
685 => 2,
686 => 3,
687 => 2,
688 => 2,
689 => 2,
690 => 2,
691 => 3,
692 => 2,
693 => 2,
694 => 3,
695 => 2,
696 => 2,
697 => 2,
698 => 2,
699 => 3,
700 => 3,
701 => 2,
702 => 2,
703 => 2,
704 => 3,
705 => 3,
706 => 3,
707 => 2,
708 => 2,
709 => 2,
710 => 2,
711 => 2,
712 => 2,
713 => 2,
714 => 2,
715 => 2,
716 => 2,
717 => 2,
718 => 2,
719 => 2,
720 => 2,
721 => 2,
722 => 3,
723 => 2,
724 => 2,
725 => 2,
726 => 3,
727 => 2,
728 => 2,
729 => 2,
730 => 2,
731 => 2,
732 => 2,
733 => 2,
734 => 2,
735 => 2,
736 => 2,
737 => 2,
738 => 2,
739 => 2,
740 => 2,
741 => 2,
742 => 2,
743 => 2,
744 => 2,
745 => 2,
746 => 2,
747 => 2,
748 => 2,
749 => 2,
750 => 2,
751 => 3,
752 => 3,
753 => 2,
754 => 2,
755 => 2,
756 => 3,
757 => 3,
758 => 3,
759 => 2,
760 => 2,
761 => 3,
762 => 2,
763 => 2,
764 => 2,
765 => 2,
766 => 2,
767 => 2,
768 => 2,
769 => 2,
770 => 3,
771 => 2,
772 => 2,
773 => 2,
774 => 2,
775 => 3,
776 => 2,
777 => 2,
778 => 3,
779 => 2,
780 => 2,
781 => 2,
782 => 2,
783 => 2,
784 => 3,
785 => 2,
786 => 3,
787 => 2,
788 => 2,
789 => 2,
790 => 2,
791 => 2,
792 => 2,
793 => 2,
794 => 2,
795 => 2,
796 => 2,
797 => 2,
798 => 2,
799 => 2,
800 => 3,
801 => 2,
802 => 2,
803 => 2,
804 => 2,
805 => 2,
806 => 2,
807 => 3,
808 => 2,
809 => 2,
810 => 2,
811 => 2,
812 => 2,
813 => 2,
814 => 2,
815 => 2,
816 => 2,
817 => 2,
818 => 2,
819 => 3,
820 => 2,
821 => 2,
822 => 2,
823 => 2,
824 => 2,
825 => 2,
826 => 2,
827 => 2,
828 => 2,
829 => 2,
830 => 2,
831 => 2,
832 => 2,
833 => 3,
834 => 2,
835 => 2,
836 => 2,
837 => 2,
838 => 2,
839 => 2,
840 => 2,
841 => 2,
842 => 2,
843 => 2,
844 => 2,
845 => 2,
846 => 2,
847 => 2,
848 => 2,
849 => 2,
850 => 2,
851 => 3,
852 => 2,
853 => 2,
854 => 2,
855 => 3,
856 => 2,
857 => 2,
858 => 2,
859 => 3,
860 => 2,
861 => 3,
862 => 3,
863 => 2,
864 => 2,
865 => 3,
866 => 3,
867 => 2,
868 => 3,
869 => 2,
870 => 2,
871 => 2,
872 => 2,
873 => 2,
874 => 2,
875 => 2,
876 => 3,
877 => 2,
878 => 2,
879 => 2,
880 => 2,
881 => 2,
882 => 2,
883 => 2,
884 => 2,
885 => 2,
886 => 2,
887 => 2,
888 => 2,
889 => 2,
890 => 2,
891 => 2,
892 => 2,
893 => 2,
894 => 2,
895 => 2,
896 => 2,
897 => 2,
898 => 2,
899 => 2,
900 => 2,
901 => 2,
902 => 2,
903 => 2,
904 => 2,
905 => 2,
906 => 2,
907 => 2,
908 => 2,
909 => 2,
910 => 2,
911 => 3,
912 => 3,
913 => 2,
914 => 2,
915 => 2,
916 => 2,
917 => 2,
918 => 2,
919 => 2,
920 => 3,
921 => 2,
922 => 2,
923 => 2,
924 => 2,
925 => 2,
926 => 2,
927 => 2,
928 => 2,
929 => 2,
930 => 2,
931 => 2,
932 => 2,
933 => 2,
934 => 2,
935 => 2,
936 => 2,
937 => 2,
938 => 2,
939 => 2,
940 => 2,
941 => 2,
942 => 2,
943 => 2,
944 => 2,
945 => 2,
946 => 3,
947 => 3,
948 => 2,
949 => 3,
950 => 3,
951 => 3,
952 => 2,
953 => 3,
954 => 2,
955 => 3,
956 => 2,
957 => 3,
958 => 2,
959 => 3,
960 => 2,
961 => 2,
962 => 3,
963 => 2,
964 => 2,
965 => 3,
966 => 3,
967 => 2,
968 => 3,
969 => 2,
970 => 2,
971 => 2,
972 => 2,
973 => 2,
974 => 2,
975 => 2,
976 => 2,
977 => 3,
978 => 3,
979 => 2,
980 => 3,
981 => 3,
982 => 2,
983 => 2,
984 => 2,
985 => 2,
986 => 2,
987 => 2,
988 => 2,
989 => 2,
990 => 3,
991 => 3,
992 => 2,
993 => 2,
994 => 2,
995 => 2,
996 => 2,
997 => 2,
998 => 2,
999 => 2,
1000 => 2,
1001 => 2,
1002 => 2,
1003 => 2,
1004 => 2,
1005 => 2,
1006 => 2,
1007 => 2,
1008 => 2,
1009 => 3,
1010 => 2,
1011 => 2,
1012 => 3,
1013 => 3,
1014 => 2,
1015 => 2,
1016 => 3,
1017 => 3,
1018 => 3,
1019 => 2,
1020 => 2,
1021 => 3,
1022 => 2,
1023 => 2,
1024 => 2,
1025 => 2,
1026 => 2,
1027 => 2,
1028 => 2,
1029 => 2,
1030 => 2,
1031 => 2,
1032 => 2,
1033 => 2,
1034 => 2,
1035 => 2,
1036 => 2,
1037 => 2,
1038 => 2,
1039 => 2,
1040 => 2,
1041 => 2,
1042 => 2,
1043 => 2,
1044 => 3,
1045 => 2,
1046 => 3,
1047 => 3,
1048 => 2,
1049 => 2,
1050 => 2,
1051 => 2,
1052 => 2,
1053 => 2,
1054 => 2,
1055 => 2,
1056 => 2,
1057 => 3,
1058 => 3,
1059 => 2,
1060 => 2,
1061 => 2,
1062 => 2,
1063 => 2,
1064 => 2,
1065 => 2,
1066 => 2,
1067 => 2,
1068 => 2,
1069 => 2,
1070 => 2,
1071 => 2,
1072 => 2,
1073 => 2,
1074 => 3,
1075 => 2,
1076 => 2,
1077 => 2,
1078 => 2,
1079 => 2,
1080 => 3,
1081 => 3,
1082 => 2,
1083 => 3,
1084 => 2,
1085 => 2,
1086 => 2,
1087 => 3,
1088 => 2,
1089 => 2,
1090 => 2,
1091 => 2,
1092 => 2,
1093 => 2,
1094 => 3,
1095 => 3,
1096 => 3,
1097 => 2,
1098 => 3,
1099 => 2,
1100 => 3,
1101 => 2,
1102 => 2,
1103 => 2,
1104 => 2,
1105 => 2,
1106 => 2,
1107 => 2,
1108 => 2,
1109 => 2,
1110 => 2,
1111 => 2,
1112 => 2,
1113 => 2,
1114 => 2,
1115 => 2,
1116 => 2,
1117 => 2,
1118 => 2,
1119 => 2,
1120 => 2,
1121 => 2,
1122 => 2,
1123 => 2,
1124 => 2,
1125 => 2,
1126 => 2,
1127 => 2,
1128 => 2,
1129 => 2,
1130 => 2,
1131 => 2,
1132 => 2,
1133 => 2,
1134 => 2,
1135 => 2,
1136 => 2,
1137 => 3,
1138 => 3,
1139 => 3,
1140 => 2,
1141 => 3,
1142 => 2,
1143 => 2,
1144 => 2,
1145 => 2,
1146 => 2,
1147 => 2,
1148 => 2,
1149 => 2,
1150 => 2,
1151 => 2,
1152 => 2,
1153 => 2,
1154 => 2,
1155 => 2,
1156 => 2,
1157 => 2,
1158 => 2,
1159 => 2,
1160 => 2,
1161 => 3,
1162 => 2,
1163 => 2,
1164 => 2,
1165 => 2,
1166 => 2,
1167 => 2,
1168 => 2,
1169 => 2,
1170 => 2,
1171 => 2,
1172 => 2,
1173 => 2,
1174 => 2,
1175 => 2,
1176 => 2,
1177 => 3,
1178 => 2,
1179 => 3,
1180 => 3,
1181 => 3,
1182 => 2,
1183 => 2,
1184 => 3,
1185 => 2,
1186 => 2,
1187 => 2,
1188 => 2,
1189 => 2,
1190 => 2,
1191 => 2,
1192 => 2,
1193 => 2,
1194 => 2,
1195 => 2,
1196 => 2,
1197 => 2,
1198 => 2,
1199 => 2,
1200 => 2,
1201 => 2,
1202 => 2,
1203 => 2,
1204 => 2,
1205 => 2,
1206 => 2,
1207 => 2,
1208 => 2,
1209 => 3,
1210 => 3,
1211 => 3,
1212 => 3,
1213 => 2,
1214 => 2,
1215 => 2,
1216 => 2,
1217 => 2,
1218 => 2,
1219 => 2,
1220 => 2,
1221 => 2,
1222 => 2,
1223 => 2,
1224 => 2,
1225 => 2,
1226 => 3,
1227 => 2,
1228 => 2,
1229 => 2,
1230 => 2,
1231 => 2,
1232 => 2,
1233 => 3,
1234 => 3,
1235 => 2,
1236 => 2,
1237 => 2,
1238 => 3,
1239 => 2,
1240 => 2,
1241 => 2,
1242 => 2,
1243 => 3,
1244 => 2,
1245 => 2,
1246 => 2,
1247 => 2,
1248 => 2,
1249 => 2,
1250 => 2,
1251 => 2,
1252 => 2,
1253 => 2,
1254 => 2,
1255 => 2,
1256 => 3,
1257 => 2,
1258 => 2,
1259 => 2,
1260 => 2,
1261 => 2,
1262 => 3,
1263 => 2,
1264 => 3,
1265 => 3,
1266 => 3,
1267 => 2,
1268 => 2,
1269 => 2,
1270 => 2,
1271 => 2,
1272 => 2,
1273 => 2,
1274 => 2,
1275 => 2,
1276 => 2,
1277 => 2,
1278 => 2,
1279 => 2,
1280 => 2,
1281 => 2,
1282 => 2,
1283 => 2,
1284 => 2,
1285 => 2,
1286 => 2,
1287 => 2,
1288 => 2,
1289 => 3,
1290 => 2,
1291 => 3,
1292 => 2,
1293 => 3,
1294 => 2,
1295 => 3,
1296 => 2,
1297 => 3,
1298 => 3,
1299 => 3,
1300 => 2,
1301 => 3,
1302 => 3,
1303 => 3,
1304 => 3,
1305 => 3,
1306 => 3,
1307 => 3,
1308 => 3,
1309 => 2,
1310 => 2,
1311 => 2,
1312 => 3,
1313 => 2,
1314 => 2,
1315 => 3,
1316 => 2,
1317 => 2,
1318 => 2,
1319 => 2,
1320 => 2,
1321 => 2,
1322 => 2,
1323 => 2,
1324 => 2,
1325 => 3,
1326 => 3,
1327 => 2,
1328 => 2,
1329 => 3,
1330 => 3,
1331 => 2,
1332 => 2,
1333 => 2,
1334 => 2,
1335 => 3,
1336 => 3,
1337 => 2,
1338 => 2,
1339 => 2,
1340 => 2,
1341 => 2,
1342 => 2,
1343 => 2,
1344 => 2,
1345 => 2,
1346 => 2,
1347 => 2,
1348 => 3,
1349 => 2,
1350 => 2,
1351 => 2,
1352 => 2,
1353 => 3,
1354 => 3,
1355 => 3,
1356 => 2,
1357 => 2,
1358 => 2,
1359 => 2,
1360 => 2,
1361 => 2,
1362 => 2,
1363 => 2,
1364 => 2,
1365 => 2,
1366 => 2,
1367 => 2,
1368 => 2,
1369 => 2,
1370 => 3,
1371 => 3,
1372 => 3,
1373 => 2,
1374 => 2,
1375 => 2,
1376 => 2,
1377 => 3,
1378 => 2,
1379 => 2,
1380 => 2,
1381 => 2,
1382 => 2,
1383 => 2,
1384 => 2,
1385 => 2,
1386 => 2,
1387 => 2,
1388 => 2,
1389 => 3,
1390 => 3,
1391 => 2,
1392 => 2,
1393 => 2,
1394 => 2,
1395 => 2,
1396 => 2,
1397 => 2,
1398 => 2,
1399 => 2,
1400 => 2,
1401 => 2,
1402 => 2,
1403 => 2,
1404 => 2,
1405 => 2,
1406 => 2,
1407 => 3,
1408 => 3,
1409 => 2,
1410 => 2,
1411 => 3,
1412 => 2,
1413 => 2,
1414 => 2,
1415 => 2,
1416 => 2,
1417 => 2,
1418 => 2,
1419 => 2,
1420 => 2,
1421 => 2,
1422 => 2,
1423 => 2,
1424 => 3,
1425 => 2,
1426 => 2,
1427 => 3,
1428 => 2,
1429 => 2,
1430 => 2,
1431 => 2,
1432 => 2,
1433 => 2,
1434 => 2,
1435 => 2,
1436 => 2,
1437 => 2,
1438 => 2,
1439 => 2,
1440 => 2,
1441 => 2,
1442 => 2,
1443 => 2,
1444 => 2,
1445 => 2,
1446 => 2,
1447 => 2,
1448 => 3,
1449 => 2,
1450 => 2,
1451 => 3,
1452 => 2,
1453 => 2,
1454 => 2,
1455 => 2,
1456 => 2,
1457 => 2,
1458 => 2,
1459 => 3,
1460 => 2,
1461 => 2,
1462 => 2,
1463 => 2,
1464 => 2,
1465 => 2,
1466 => 2,
1467 => 2,
1468 => 3,
1469 => 3,
1470 => 3,
1471 => 2,
1472 => 3,
1473 => 2,
1474 => 2,
1475 => 2,
1476 => 2,
1477 => 2,
1478 => 2,
1479 => 2,
1480 => 2,
1481 => 2,
1482 => 3,
1483 => 3,
1484 => 3,
1485 => 3,
1486 => 2,
1487 => 3,
1488 => 3,
1489 => 3,
1490 => 3,
1491 => 3,
1492 => 2,
1493 => 3,
1494 => 2,
1495 => 2,
1496 => 3,
1497 => 3,
1498 => 2,
1499 => 2,
1500 => 3,
1501 => 2,
1502 => 3,
1503 => 3,
1504 => 3,
1505 => 3,
1506 => 2,
1507 => 2,
1508 => 2,
1509 => 2,
1510 => 3,
1511 => 3,
1512 => 2,
1513 => 3,
1514 => 2,
1515 => 3,
1516 => 2,
1517 => 2,
1518 => 2,
1519 => 2,
1520 => 3,
1521 => 3,
1522 => 2,
1523 => 2,
1524 => 2,
1525 => 2,
1526 => 2,
1527 => 2,
1528 => 2,
1529 => 2,
1530 => 3,
1531 => 2,
1532 => 2,
1533 => 2,
1534 => 2,
1535 => 2,
1536 => 2,
1537 => 2,
1538 => 2,
1539 => 2,
1540 => 2,
1541 => 2,
1542 => 3,
1543 => 2,
1544 => 2,
1545 => 2,
1546 => 2,
1547 => 2,
1548 => 3,
1549 => 2,
1550 => 2,
1551 => 2,
1552 => 2,
1553 => 2,
1554 => 2,
1555 => 2,
1556 => 3,
1557 => 2,
1558 => 2,
1559 => 2,
1560 => 2,
1561 => 2,
1562 => 2,
1563 => 2,
1564 => 2,
1565 => 3,
1566 => 3,
1567 => 2,
1568 => 2,
1569 => 2,
1570 => 2,
1571 => 3,
1572 => 2,
1573 => 2,
1574 => 2,
1575 => 2,
1576 => 3,
1577 => 3,
1578 => 2,
1579 => 2,
1580 => 2,
1581 => 2,
1582 => 2,
1583 => 3,
1584 => 2,
1585 => 2,
1586 => 2,
1587 => 2,
1588 => 2,
1589 => 2,
1590 => 2,
1591 => 2,
1592 => 2,
1593 => 2,
1594 => 2,
1595 => 2,
1596 => 3,
1597 => 2,
1598 => 2,
1599 => 2,
1600 => 2,
1601 => 2,
1602 => 2,
1603 => 2,
1604 => 2,
1605 => 3,
1606 => 2,
1607 => 3,
1608 => 2,
1609 => 2,
1610 => 3,
1611 => 2,
1612 => 3,
1613 => 2,
1614 => 2,
1615 => 2,
1616 => 2,
1617 => 2,
1618 => 2,
1619 => 2,
1620 => 2,
1621 => 2,
1622 => 2,
1623 => 2,
1624 => 2,
1625 => 2,
1626 => 2,
1627 => 2,
1628 => 2,
1629 => 2,
1630 => 2,
1631 => 2,
1632 => 2,
1633 => 2,
1634 => 2,
1635 => 2,
1636 => 2,
1637 => 2,
1638 => 2,
1639 => 2,
1640 => 2,
1641 => 2,
1642 => 2,
1643 => 2,
1644 => 2,
1645 => 2,
1646 => 2,
1647 => 2,
1648 => 3,
1649 => 2,
1650 => 2,
1651 => 3,
1652 => 3,
1653 => 3,
1654 => 2,
1655 => 2,
1656 => 2,
1657 => 3,
1658 => 3,
1659 => 2,
1660 => 3,
1661 => 2,
1662 => 2,
1663 => 2,
1664 => 2,
1665 => 2,
1666 => 2,
1667 => 2,
1668 => 3,
1669 => 3,
1670 => 2,
1671 => 2,
1672 => 2,
1673 => 2,
1674 => 2,
1675 => 2,
1676 => 2,
1677 => 3,
1678 => 2,
1679 => 2,
1680 => 3,
1681 => 2,
1682 => 2,
1683 => 3,
1684 => 3,
1685 => 3,
1686 => 2,
1687 => 2,
1688 => 2,
1689 => 2,
1690 => 2,
1691 => 2,
1692 => 2,
1693 => 2,
1694 => 2,
1695 => 2,
1696 => 2,
1697 => 2,
1698 => 2,
1699 => 2,
1700 => 2,
1701 => 2,
1702 => 3,
1703 => 2,
1704 => 2,
1705 => 2,
1706 => 2,
1707 => 2,
1708 => 2,
1709 => 2,
1710 => 2,
1711 => 2,
1712 => 2,
1713 => 3,
1714 => 2,
1715 => 2,
1716 => 2,
1717 => 2,
1718 => 2,
1719 => 2,
1720 => 3,
1721 => 2,
1722 => 2,
1723 => 2,
1724 => 2,
1725 => 2,
1726 => 3,
1727 => 2,
1728 => 2,
1729 => 2,
1730 => 2,
1731 => 2,
1732 => 2,
1733 => 2,
1734 => 2,
1735 => 2,
1736 => 2,
1737 => 2,
1738 => 2,
1739 => 2,
1740 => 2,
1741 => 2,
1742 => 2,
1743 => 2,
1744 => 2,
1745 => 2,
1746 => 2,
1747 => 2,
1748 => 2,
1749 => 2,
1750 => 2,
1751 => 3,
1752 => 2,
1753 => 2,
1754 => 2,
1755 => 2,
1756 => 2,
1757 => 2,
1758 => 2,
1759 => 2,
1760 => 2,
1761 => 2,
1762 => 2,
1763 => 3,
1764 => 3,
1765 => 2,
1766 => 3,
1767 => 2,
1768 => 3,
1769 => 3,
1770 => 2,
1771 => 2,
1772 => 2,
1773 => 2,
1774 => 2,
1775 => 2,
1776 => 2,
1777 => 2,
1778 => 2,
1779 => 2,
1780 => 2,
1781 => 2,
1782 => 2,
1783 => 2,
1784 => 2,
1785 => 2,
1786 => 3,
1787 => 2,
1788 => 2,
1789 => 3,
1790 => 2,
1791 => 3,
1792 => 2,
1793 => 2,
1794 => 2,
1795 => 2,
1796 => 2,
1797 => 2,
1798 => 2,
1799 => 2,
1800 => 3,
1801 => 2,
1802 => 2,
1803 => 2,
1804 => 2,
1805 => 3,
1806 => 2,
1807 => 2,
1808 => 2,
1809 => 2,
1810 => 3,
1811 => 2,
1812 => 2,
1813 => 3,
1814 => 2,
1815 => 2,
1816 => 3,
1817 => 2,
1818 => 2,
1819 => 2,
1820 => 3,
1821 => 3,
1822 => 2,
1823 => 2,
1824 => 2,
1825 => 2,
1826 => 2,
1827 => 2,
1828 => 2,
1829 => 2,
1830 => 3,
1831 => 2,
1832 => 2,
1833 => 3,
1834 => 2,
1835 => 2,
1836 => 2,
1837 => 3,
1838 => 3,
1839 => 2,
1840 => 3,
1841 => 3,
1842 => 2,
1843 => 2,
1844 => 2,
1845 => 2,
1846 => 2,
1847 => 2,
1848 => 2,
1849 => 2,
1850 => 2,
1851 => 2,
1852 => 2,
1853 => 2,
1854 => 2,
1855 => 2,
1856 => 2,
1857 => 2,
1858 => 2,
1859 => 2,
1860 => 2,
1861 => 2,
1862 => 3,
1863 => 2,
1864 => 2,
1865 => 2,
1866 => 2,
1867 => 2,
1868 => 2,
1869 => 2,
1870 => 2,
1871 => 2,
1872 => 2,
1873 => 2,
1874 => 3,
1875 => 2,
1876 => 2,
1877 => 2,
1878 => 2,
1879 => 2,
1880 => 3,
1881 => 2,
1882 => 2,
1883 => 3,
1884 => 3,
1885 => 2,
1886 => 2,
1887 => 2,
1888 => 2,
1889 => 2,
1890 => 2,
1891 => 2,
1892 => 3,
1893 => 3,
1894 => 2,
1895 => 2,
1896 => 2,
1897 => 2,
1898 => 2,
1899 => 2,
1900 => 3,
1901 => 3,
1902 => 2,
1903 => 2,
1904 => 2,
1905 => 2,
1906 => 2,
1907 => 2,
1908 => 2,
1909 => 2,
1910 => 2,
1911 => 2,
1912 => 2,
1913 => 3,
1914 => 3,
1915 => 3,
1916 => 2,
1917 => 3,
1918 => 2,
1919 => 2,
1920 => 2,
1921 => 2,
1922 => 2,
1923 => 2,
1924 => 2,
1925 => 2,
1926 => 2,
1927 => 2,
1928 => 2,
1929 => 2,
1930 => 2,
1931 => 2,
1932 => 2,
1933 => 2,
1934 => 2,
1935 => 2,
1936 => 2,
1937 => 2,
1938 => 2,
1939 => 2,
1940 => 3,
1941 => 2,
1942 => 2,
1943 => 2,
1944 => 2,
1945 => 2,
1946 => 3,
1947 => 3,
1948 => 2,
1949 => 3,
1950 => 3,
1951 => 3,
1952 => 2,
1953 => 2,
1954 => 2,
1955 => 2,
1956 => 3,
1957 => 2,
1958 => 3,
1959 => 2,
1960 => 2,
1961 => 2,
1962 => 2,
1963 => 3,
1964 => 2,
1965 => 2,
1966 => 2,
1967 => 3,
1968 => 2,
1969 => 2,
1970 => 2,
1971 => 2,
1972 => 2,
1973 => 2,
1974 => 2,
1975 => 2,
1976 => 2,
1977 => 2,
1978 => 3,
1979 => 2,
1980 => 2,
1981 => 2,
1982 => 2,
1983 => 2,
1984 => 2,
1985 => 3,
1986 => 2,
1987 => 2,
1988 => 2,
1989 => 2,
1990 => 2,
1991 => 2,
1992 => 3,
1993 => 2,
1994 => 2,
1995 => 2,
1996 => 2,
1997 => 2,
1998 => 2,
1999 => 2,
2000 => 2,
2001 => 2,
2002 => 2,
2003 => 3,
2004 => 3,
2005 => 3,
2006 => 2,
2007 => 2,
2008 => 2,
2009 => 3,
2010 => 2,
2011 => 2,
2012 => 2,
2013 => 2,
2014 => 2,
2015 => 3,
2016 => 2,
2017 => 3,
2018 => 2,
2019 => 3,
2020 => 3,
2021 => 3,
2022 => 2,
2023 => 2,
2024 => 2,
2025 => 3,
2026 => 2,
2027 => 2,
2028 => 2,
2029 => 2,
2030 => 2,
2031 => 2,
2032 => 2,
2033 => 2,
2034 => 2,
2035 => 2,
2036 => 3,
2037 => 2,
2038 => 2,
2039 => 3,
2040 => 3,
2041 => 3,
2042 => 3,
2043 => 2,
2044 => 2,
2045 => 2,
2046 => 3,
2047 => 3,
2048 => 2,
2049 => 2,
2050 => 2,
2051 => 2,
2052 => 2,
2053 => 2,
2054 => 2,
2055 => 2,
2056 => 2,
2057 => 2,
2058 => 2,
2059 => 2,
2060 => 2,
2061 => 3,
2062 => 2,
2063 => 2,
2064 => 2,
2065 => 2,
2066 => 2,
2067 => 3,
2068 => 2,
2069 => 2,
2070 => 3,
2071 => 2,
2072 => 3,
2073 => 3,
2074 => 3,
2075 => 2,
2076 => 3,
2077 => 2,
2078 => 2,
2079 => 2,
2080 => 2,
2081 => 2,
2082 => 2,
2083 => 2,
2084 => 3,
2085 => 2,
2086 => 2,
2087 => 2,
2088 => 2,
2089 => 3,
2090 => 3,
2091 => 3,
2092 => 3,
2093 => 2,
2094 => 2,
2095 => 3,
2096 => 3,
2097 => 2,
2098 => 2,
2099 => 2,
2100 => 2,
2101 => 2,
2102 => 3,
2103 => 3,
2104 => 3,
2105 => 3,
2106 => 3,
2107 => 2,
2108 => 2,
2109 => 2,
2110 => 2,
2111 => 2,
2112 => 2,
2113 => 2,
2114 => 2,
2115 => 2,
2116 => 2,
2117 => 2,
2118 => 2,
2119 => 2,
2120 => 2,
2121 => 2,
2122 => 2,
2123 => 2,
2124 => 2,
2125 => 2,
2126 => 2,
2127 => 2,
2128 => 2,
2129 => 2,
2130 => 2,
2131 => 2,
2132 => 2,
2133 => 2,
2134 => 2,
2135 => 2,
2136 => 2,
2137 => 2,
2138 => 2,
2139 => 2,
2140 => 2,
2141 => 2,
2142 => 3,
2143 => 2,
2144 => 2,
2145 => 2,
2146 => 3,
2147 => 2,
2148 => 2,
2149 => 2,
2150 => 2,
2151 => 2,
2152 => 2,
2153 => 3,
2154 => 2,
2155 => 2,
2156 => 2,
2157 => 2,
2158 => 2,
2159 => 2,
2160 => 2,
2161 => 2,
2162 => 2,
2163 => 2,
2164 => 3,
2165 => 3,
2166 => 3,
2167 => 3,
2168 => 2,
2169 => 2,
2170 => 3,
2171 => 2,
2172 => 2,
2173 => 2,
2174 => 3,
2175 => 2,
2176 => 2,
2177 => 2,
2178 => 2,
2179 => 2,
2180 => 2,
2181 => 3,
2182 => 2,
2183 => 2,
2184 => 2,
2185 => 2,
2186 => 3,
2187 => 2,
2188 => 2,
2189 => 3,
2190 => 2,
2191 => 2,
2192 => 3,
2193 => 2,
2194 => 2,
2195 => 2,
2196 => 2,
2197 => 3,
2198 => 2,
2199 => 3,
2200 => 2,
2201 => 2,
2202 => 2,
2203 => 2,
2204 => 3,
2205 => 3,
2206 => 3,
2207 => 2,
2208 => 2,
2209 => 2,
2210 => 2,
2211 => 2,
2212 => 2,
2213 => 2,
2214 => 2,
2215 => 2,
2216 => 2,
2217 => 2,
2218 => 2,
2219 => 2,
2220 => 2,
2221 => 2,
2222 => 2,
2223 => 2,
2224 => 2,
2225 => 2,
2226 => 2,
2227 => 2,
2228 => 2,
2229 => 2,
2230 => 3,
2231 => 2,
2232 => 2,
2233 => 2,
2234 => 2,
2235 => 2,
2236 => 2,
2237 => 2,
2238 => 3,
2239 => 2,
2240 => 2,
2241 => 2,
2242 => 2,
2243 => 2,
2244 => 2,
2245 => 3,
2246 => 2,
2247 => 2,
2248 => 2,
2249 => 2,
2250 => 2,
2251 => 2,
2252 => 3,
2253 => 3,
2254 => 2,
2255 => 2,
2256 => 2,
2257 => 2,
2258 => 2,
2259 => 2,
2260 => 2,
2261 => 2,
2262 => 2,
2263 => 2,
2264 => 3,
2265 => 3,
2266 => 2,
2267 => 2,
2268 => 2,
2269 => 2,
2270 => 2,
2271 => 2,
2272 => 2,
2273 => 3,
2274 => 2,
2275 => 3,
2276 => 2,
2277 => 2,
2278 => 3,
2279 => 3,
2280 => 2,
2281 => 2,
2282 => 2,
2283 => 2,
2284 => 2,
2285 => 2,
2286 => 2,
2287 => 3,
2288 => 2,
2289 => 3,
2290 => 3,
2291 => 3,
2292 => 3,
2293 => 2,
2294 => 2,
2295 => 2,
2296 => 2,
2297 => 2,
2298 => 2,
2299 => 2,
2300 => 2,
2301 => 2,
2302 => 2,
2303 => 2,
2304 => 2,
2305 => 2,
2306 => 2,
2307 => 2,
2308 => 2,
2309 => 2,
2310 => 2,
2311 => 2,
2312 => 2,
2313 => 2,
2314 => 2,
2315 => 2,
2316 => 2,
2317 => 2,
2318 => 3,
2319 => 2,
2320 => 3,
2321 => 3,
2322 => 3,
2323 => 2,
2324 => 2,
2325 => 2,
2326 => 2,
2327 => 2,
2328 => 2,
2329 => 3,
2330 => 2,
2331 => 2,
2332 => 2,
2333 => 2,
2334 => 2,
2335 => 2,
2336 => 2,
2337 => 3,
2338 => 3,
2339 => 3,
2340 => 2,
2341 => 3,
2342 => 2,
2343 => 2,
2344 => 2,
2345 => 2,
2346 => 3,
2347 => 3,
2348 => 2,
2349 => 2,
2350 => 3,
2351 => 3,
2352 => 2,
2353 => 2,
2354 => 3,
2355 => 2,
2356 => 3,
2357 => 2,
2358 => 2,
2359 => 2,
2360 => 2,
2361 => 2,
2362 => 2,
2363 => 2,
2364 => 2,
2365 => 3,
2366 => 2,
2367 => 2,
2368 => 3,
2369 => 3,
2370 => 2,
2371 => 2,
2372 => 2,
2373 => 2,
2374 => 3,
2375 => 2,
2376 => 2,
2377 => 2,
2378 => 3,
2379 => 2,
2380 => 2,
2381 => 2,
2382 => 3,
2383 => 3,
2384 => 2,
2385 => 2,
2386 => 3,
2387 => 2,
2388 => 2,
2389 => 2,
2390 => 2,
2391 => 2,
2392 => 2,
2393 => 2,
2394 => 2,
2395 => 3,
2396 => 2,
2397 => 2,
2398 => 2,
2399 => 2,
2400 => 2,
2401 => 2,
2402 => 2,
2403 => 2,
2404 => 2,
2405 => 2,
2406 => 2,
2407 => 2,
2408 => 2,
2409 => 2,
2410 => 2,
2411 => 2,
2412 => 3,
2413 => 2,
2414 => 2,
2415 => 2,
2416 => 2,
2417 => 2,
2418 => 2,
2419 => 2,
2420 => 2,
2421 => 2,
2422 => 2,
2423 => 2,
2424 => 2,
2425 => 3,
2426 => 2,
2427 => 2,
2428 => 3,
2429 => 3,
2430 => 2,
2431 => 2,
2432 => 2,
2433 => 3,
2434 => 2,
2435 => 2,
2436 => 3,
2437 => 3,
2438 => 3,
2439 => 2,
2440 => 2,
2441 => 3,
2442 => 2,
2443 => 2,
2444 => 2,
2445 => 3,
2446 => 2,
2447 => 2,
2448 => 3,
2449 => 2,
2450 => 2,
2451 => 2,
2452 => 2,
2453 => 2,
2454 => 2,
2455 => 2,
2456 => 3,
2457 => 3,
2458 => 2,
2459 => 2,
2460 => 3,
2461 => 2,
2462 => 2,
2463 => 3,
2464 => 2,
2465 => 2,
2466 => 2,
2467 => 2,
2468 => 2,
2469 => 2,
2470 => 2,
2471 => 2,
2472 => 2,
2473 => 2,
2474 => 2,
2475 => 2,
2476 => 2,
2477 => 2,
2478 => 2,
2479 => 3,
2480 => 2,
2481 => 2,
2482 => 2,
2483 => 2,
2484 => 2,
2485 => 3,
2486 => 2,
2487 => 2,
2488 => 2,
2489 => 2,
2490 => 3,
2491 => 3,
2492 => 3,
2493 => 3,
2494 => 2,
2495 => 2,
2496 => 3,
2497 => 2,
2498 => 2,
2499 => 2,
2500 => 2,
2501 => 3,
2502 => 2,
2503 => 2,
2504 => 2,
2505 => 2,
2506 => 2,
2507 => 2,
2508 => 2,
2509 => 2,
2510 => 3,
2511 => 3,
2512 => 2,
2513 => 3,
2514 => 2,
2515 => 2,
2516 => 2,
2517 => 2,
2518 => 2,
2519 => 2,
2520 => 2,
2521 => 2,
2522 => 2,
2523 => 2,
2524 => 2,
2525 => 2,
2526 => 2,
2527 => 2,
2528 => 2,
2529 => 2,
2530 => 2,
2531 => 2,
2532 => 2,
2533 => 2,
2534 => 2,
2535 => 3,
2536 => 3,
2537 => 3,
2538 => 2,
2539 => 3,
2540 => 3,
2541 => 2,
2542 => 3,
2543 => 3,
2544 => 3,
2545 => 2,
2546 => 2,
2547 => 2,
2548 => 2,
2549 => 2,
2550 => 2,
2551 => 2,
2552 => 2,
2553 => 3,
2554 => 2,
2555 => 3,
2556 => 2,
2557 => 2,
2558 => 2,
2559 => 2,
2560 => 2,
2561 => 2,
2562 => 2,
2563 => 2,
2564 => 2,
2565 => 2,
2566 => 2,
2567 => 2,
2568 => 3,
2569 => 2,
2570 => 2,
2571 => 2,
2572 => 2,
2573 => 2,
2574 => 2,
2575 => 2,
2576 => 2,
2577 => 2,
2578 => 2,
2579 => 2,
2580 => 3,
2581 => 3,
2582 => 3,
2583 => 3,
2584 => 3,
2585 => 2,
2586 => 2,
2587 => 3,
2588 => 2,
2589 => 3,
2590 => 3,
2591 => 2,
2592 => 3,
2593 => 2,
2594 => 2,
2595 => 3,
2596 => 2,
2597 => 3,
2598 => 3,
2599 => 2,
2600 => 2,
2601 => 2,
2602 => 2,
2603 => 2,
2604 => 2,
2605 => 2,
2606 => 2,
2607 => 2,
2608 => 3,
2609 => 2,
2610 => 2,
2611 => 3,
2612 => 3,
2613 => 2,
2614 => 2,
2615 => 2,
2616 => 3,
2617 => 2,
2618 => 2,
2619 => 2,
2620 => 2,
2621 => 2,
2622 => 2,
2623 => 2,
2624 => 2,
2625 => 2,
2626 => 3,
2627 => 2,
2628 => 2,
2629 => 2,
2630 => 2,
2631 => 2,
2632 => 2,
2633 => 2,
2634 => 2,
2635 => 2,
2636 => 2,
2637 => 2,
2638 => 2,
2639 => 2,
2640 => 2,
2641 => 3,
2642 => 3,
2643 => 2,
2644 => 2,
2645 => 3,
2646 => 3,
2647 => 2,
2648 => 3,
2649 => 2,
2650 => 2,
2651 => 2,
2652 => 2,
2653 => 3,
2654 => 2,
2655 => 2,
2656 => 3,
2657 => 2,
2658 => 2,
2659 => 2,
2660 => 2,
2661 => 2,
2662 => 2,
2663 => 2,
2664 => 2,
2665 => 2,
2666 => 2,
2667 => 2,
2668 => 2,
2669 => 2,
2670 => 3,
2671 => 3,
2672 => 2,
2673 => 2,
2674 => 3,
2675 => 3,
2676 => 2,
2677 => 2,
2678 => 2,
2679 => 3,
2680 => 2,
2681 => 2,
2682 => 2,
2683 => 2,
2684 => 2,
2685 => 2,
2686 => 2,
2687 => 2,
2688 => 2,
2689 => 2,
2690 => 2,
2691 => 2,
2692 => 2,
2693 => 2,
2694 => 2,
2695 => 2,
2696 => 2,
2697 => 2,
2698 => 2,
2699 => 2,
2700 => 2,
2701 => 2,
2702 => 2,
2703 => 2,
2704 => 2,
2705 => 2,
2706 => 3,
2707 => 3,
2708 => 2,
2709 => 2,
2710 => 2,
2711 => 3,
2712 => 2,
2713 => 2,
2714 => 2,
2715 => 2,
2716 => 2,
2717 => 2,
2718 => 3,
2719 => 2,
2720 => 2,
2721 => 2,
2722 => 2,
2723 => 3,
2724 => 2,
2725 => 2,
2726 => 2,
2727 => 2,
2728 => 3,
2729 => 2,
2730 => 2,
2731 => 2,
2732 => 2,
2733 => 2,
2734 => 2,
2735 => 2,
2736 => 2,
2737 => 2,
2738 => 2,
2739 => 2,
2740 => 2,
2741 => 2,
2742 => 2,
2743 => 2,
2744 => 2,
2745 => 2,
2746 => 2,
2747 => 2,
2748 => 2,
2749 => 2,
2750 => 2,
2751 => 2,
2752 => 2,
2753 => 2,
2754 => 2,
2755 => 2,
2756 => 2,
2757 => 3,
2758 => 2,
2759 => 3,
2760 => 2,
2761 => 2,
2762 => 2,
2763 => 2,
2764 => 2,
2765 => 2,
2766 => 2,
2767 => 2,
2768 => 2,
2769 => 3,
2770 => 3,
2771 => 3,
2772 => 2,
2773 => 2,
2774 => 3,
2775 => 2,
2776 => 3,
2777 => 3,
2778 => 3,
2779 => 3,
2780 => 2,
2781 => 2,
2782 => 2,
2783 => 2,
2784 => 2,
2785 => 2,
2786 => 3,
2787 => 2,
2788 => 2,
2789 => 2,
2790 => 2,
2791 => 2,
2792 => 2,
2793 => 2,
2794 => 3,
2795 => 3,
2796 => 2,
2797 => 3,
2798 => 3,
2799 => 3,
2800 => 3,
2801 => 3,
2802 => 2,
2803 => 2,
2804 => 2,
2805 => 2,
2806 => 2,
2807 => 2,
2808 => 2,
2809 => 2,
2810 => 2,
2811 => 2,
2812 => 2,
2813 => 2,
2814 => 2,
2815 => 2,
2816 => 3,
2817 => 3,
2818 => 2,
2819 => 2,
2820 => 2,
2821 => 2,
2822 => 2,
2823 => 2,
2824 => 2,
2825 => 2,
2826 => 3,
2827 => 2,
2828 => 2,
2829 => 2,
2830 => 2,
2831 => 2,
2832 => 3,
2833 => 2,
2834 => 2,
2835 => 2,
2836 => 2,
2837 => 2,
2838 => 3,
2839 => 2,
2840 => 2,
2841 => 2,
2842 => 2,
2843 => 2,
2844 => 2,
2845 => 2,
2846 => 3,
2847 => 2,
2848 => 2,
2849 => 2,
2850 => 2,
2851 => 3,
2852 => 2,
2853 => 2,
2854 => 2,
2855 => 2,
2856 => 2,
2857 => 3,
2858 => 3,
2859 => 2,
2860 => 2,
2861 => 2,
2862 => 2,
2863 => 2,
2864 => 2,
2865 => 2,
2866 => 3,
2867 => 2,
2868 => 2,
2869 => 2,
2870 => 2,
2871 => 2,
2872 => 2,
2873 => 2,
2874 => 2,
2875 => 3,
2876 => 3,
2877 => 3,
2878 => 3,
2879 => 3,
2880 => 3,
2881 => 3,
2882 => 3,
2883 => 3,
2884 => 2,
2885 => 2,
2886 => 2,
2887 => 2,
2888 => 2,
2889 => 2,
2890 => 2,
2891 => 2,
2892 => 2,
2893 => 2,
2894 => 3,
2895 => 3,
2896 => 2,
2897 => 2,
2898 => 3,
2899 => 3,
2900 => 2,
2901 => 3,
2902 => 2,
2903 => 2,
2904 => 2,
2905 => 2,
2906 => 2,
2907 => 2,
2908 => 2,
2909 => 2,
2910 => 2,
2911 => 2,
2912 => 3);

constant Nstage : integer := 25;

--constant SE : integer :=
--constant SV : integer :=
--constant FE : integer :=
--constant FV : integer :=
--constant GTE: integer :=
--constant GTV: integer :=
--constant LSE: integer :=
--constant LSV: integer :=
type Mean is array (0 to 3) of integer;
type Var is array (0 to 3) of integer;
type R is array (0 to 3) of integer;

type Rectangle is
record 
	x	: integer;
	y	: integer;
	h	: integer;
	w	: integer;
	weight : integer;
end record;

type Rectangles is array (0 to 2) of Rectangle;
type R_tab is array (0 to 2) of R;


type Feature is 
record
	--rects 		: Rectangles;
	threshold	: integer;
	nr				: integer; -- number of rectangles per feature
	greater		: integer;
	lower 		: integer; 
	ad_rectangle : integer;
end record;

--type Features is array (0 to 37) of Feature; --useless

--type Stage is
--record
	--feats			: Features;
	--threshold	: integer;
	--nf				: integer; --number of features per stage
--end record; 

type Stage is
record
	threshold : integer;
	ad_feature: integer;
	nf : integer;
end record;

type Detector is
record
	x	: integer;
	y 	: integer;
end record;

--function StageEval (signal d: in Detector; signal stageAdress : in unsigned (5 downto 0)) return integer;  
function FeatureEval(signal r_tab: in R_tab; signal rect: in Rectangles) return integer;
function test_Feature( signal sumf_q : in integer; signal meanP : in Mean; signal varP : in Var; calcul : integer; signal f_q : in Feature) return boolean;

-- procedure <procedure_name> (<type_declaration> <constant_name>	: in <type_declaration>);
--

end FACE_DETECTION_PCK;

package body FACE_DETECTION_PCK is

function StageEval (signal d: in Detector; signal stageAdress : in unsigned (5 downto 0)) return integer is
begin
	--todo
	return 0;
end;

function FeatureEval(signal r_tab : in R_tab; signal rect : in Rectangles) return integer is
variable cont1 : integer;
variable cont2 : integer;
variable cont3 : integer;
variable sum: integer;

begin
	cont1 := r_tab(0)(3)+r_tab(0)(1)-r_tab(0)(2)-r_tab(0)(3);
	cont2 := r_tab(1)(3)+r_tab(1)(1)-r_tab(1)(2)-r_tab(1)(3);
	cont3 := r_tab(2)(3)+r_tab(2)(1)-r_tab(2)(2)-r_tab(2)(3);
	
	sum := cont1*rect(0).weight + cont2*rect(1).weight + cont3*rect(2).weight;
	
	return sum;
end;


function test_Feature( signal sumf_q : in integer; signal meanP : in Mean; signal varP : in Var; calcul : integer; signal f_q : in Feature) return boolean is
variable mean : integer;
variable sq_mean : integer;
variable var_sq : integer;
variable seuil : integer;
begin
mean := meanP(4)+meanP(1)-meanP(2)-meanP(3);
sq_mean := varP(4)+varP(1)-varP(2)-varP(3);
var_sq := sq_mean*24*24-mean*mean;

seuil:= f_q.threshold;
if(sumf_q*sumf_q>=seuil*seuil*var_sq) then
	return true;
else
	return false;
end if;
end;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;


end FACE_DETECTION_PCK;