----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:49:01 06/05/2015 
-- Design Name: 
-- Module Name:    RAM_Classifier - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


--Stages--
entity ram_Stages is
port ( 	clk : in std_logic;
			adress : in integer;
			data_o : out unsigned(27 downto 0)
     );
end ram_Stages;

architecture Behavioral of ram_Stages is



type ram_t is array (0 to 24) of unsigned(27 downto 0);
signal ram : ram_t := 
(
0 => "0000000000001011000000000000",
1 => "0000000000000011000000001001",
2 => "0000000000000011000000011001",
3 => "0000000000000011000000110100",
4 => "0000000000000011000001010100",
5 => "0000000000000011000010001000",
6 => "0000000000000011000010111101",
7 => "0000000001100001000011111011",
8 => "1100001010000101000101000011",
9 => "0000000001100011000110010110",
10 => "1100001000010100000111110001",
11 => "1100010010001010001001010100",
12 => "0000000000011001001011000111",
13 => "0000000011000101001101000110",
14 => "0000110010010011001111001101",
15 => "0000000000011001010001010101",
16 => "0000000000011001010011011110",
17 => "0000000001100101010101111101",
18 => "0000000000001101011000011000",
19 => "0000000000001101011011000001",
20 => "0000000000110011011110000101",
21 => "0000000011001011100001001010",
22 => "0000000000110011100011111111",
23 => "0011001010000101100111000110",
24 => "0000011010000001101010011001"
);
begin

--process for read and write operation.
PROCESS(clk)
BEGIN
    if(rising_edge(clk)) then
        data_o <= ram(adress);
    end if;
END PROCESS;

end Behavioral;



library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

--Features--

entity ram_Features is
port ( 	clk : in std_logic;
			adress : in integer;
			data_o : out unsigned(60 downto 0)
     );
end ram_Features;

architecture Behavioral of ram_Features is

--Declaration of type and signal of a 256 element RAM
--with each element being 8 bit wide.
type ram_t is array (0 to 2912) of unsigned(60 downto 0);
signal ram : ram_t := 
(
0 => "0000000000000001000000000100001100000000000000110000000000000",
1 => "0000000000000001000000000000001100000000010101010000000000010",
2 => "0000000000000011000000000000001100000100010000000000000000100",
3 => "0000000000000011000000000000001100000000000100110000000000110",
4 => "0000000000000001000000000000001100000001010000110000000001000",
5 => "0000000000000001000000000000100100000000000000110000000001010",
6 => "0000000000000011000000000000001100000000000000010000000001100",
7 => "0000000000000001000000000000001100000000000000010000000001110",
8 => "0000000000000001000000000000001100000000000000010000000010000",
9 => "0000000000000001000000000000010100000000000000110000000010010",
10 => "0000000000010101000000000000001100000000000100110000000010100",
11 => "0000000000001011000000000000001100000000000000110000000010110",
12 => "0000000000000011000000000000001100000000000000010000000011000",
13 => "0000010010100101000000010001001000000000000000110000000011010",
14 => "0000000000000001000000000000001100000000000000010000000011100",
15 => "0000000000010001000000000000001100000010001001000000000011110",
16 => "0000000000010011000000000000001100000000000000010000000100000",
17 => "0000000000000001000000000000000100000000000000110000000100010",
18 => "0000000000000001000000100101000100000000000000110000000100100",
19 => "0000000001000001000000000000001100000000000010110000000100110",
20 => "0000000000000001000000000000001100000000000000110000000101000",
21 => "0000000000000001000000000000100100000000000000110000000101010",
22 => "0000000000000001000000000000001100000001001001010000000101100",
23 => "0000000000010101000000000000001100000000000000010000000101110",
24 => "0000000000000011000000000000000100000000000000110000000110000",
25 => "0000000000001001000000000000001100000000000000110000000110010",
26 => "0000010000001000000000000000001100000100000000000000000110100",
27 => "0000000000000001000000000000000100000000000000110000000110110",
28 => "0000000000000001000000000000001100000000000000010000000111000",
29 => "0000000000000001000000000000001100000000000000010000000111010",
30 => "0000000000010001000000000000001100000000000100010000000111100",
31 => "0000000000000001000000000000001100000000000000110000000111110",
32 => "0000000000000001000000000000001100000000000000110000001000000",
33 => "0000000000000001000000000000001100000000000001010000001000010",
34 => "0000000000000001000000000001000100000000000000110000001000100",
35 => "0000000000000001000000000000001100000000000001010000001000110",
36 => "0000000000001011000000010010001000000000000000110000001001001",
37 => "0000000000000001000000000000001100000000000000010000001001011",
38 => "0000000000000001000000000000001100000000001010010000001001101",
39 => "0000000000000001000000000000000100000000000000110000001001111",
40 => "0000000000000001000000000000000100000000000000110000001010001",
41 => "0000000000000011000000000000001100000000000000010000001010011",
42 => "0000000000000101000000000000001100000000000000010000001010101",
43 => "0000000000001001000000000000001100000000000000010000001010111",
44 => "0000010100010010000000000000101100000000000000110000001011001",
45 => "0000000000000001000000000000000100000000000000110000001011011",
46 => "0000000000000001000000000000001100000000000000010000001011101",
47 => "0000000000000001000000000001000100000000000000110000001011111",
48 => "0000000000000001000000000000001100000000010010010000001100001",
49 => "0000000001000101000000000000001100000000000000010000001100100",
50 => "0000000000000001000000000000001100000000010001010000001100110",
51 => "0000000000000001000000000000001100000000000000010000001101000",
52 => "0000000000000001000000000010010100000000000000110000001101010",
53 => "0000000001000001000000000000001100000000000000010000001101100",
54 => "0000001001010101000000000000001100000000000000110000001101110",
55 => "0000000000000001000000000000001100000010000100000000001110000",
56 => "0000000000000001000000000000001100000000010010110000001110010",
57 => "0000000000010011000000000000001100000000010010110000001110101",
58 => "0000000000101001000000000000001100000000000000010000001110111",
59 => "0000000000000111000000000000001100000000000000110000001111001",
60 => "0000000000010011000000000000001100000000000010010000001111011",
61 => "0000000000000001000000000000001100000000000000010000001111101",
62 => "0000000000010011000000000000001100000000000000110000001111111",
63 => "0000000000000001000000000000000100000000000000110000010000010",
64 => "0000000010001011000000000000001100000000000000110000010000100",
65 => "0000000000000001000000000000001100000000000000110000010000110",
66 => "0000000000000001000000000000000100000000000000110000010001000",
67 => "0000000000000001000000000000001100000000000000010000010001010",
68 => "0000000000000001000000000000001100000000000000110000010001100",
69 => "0000000000000001000000000000001100000000010100010000010001110",
70 => "0000000000000001000000000000001100000000000000010000010010000",
71 => "0000000000000011000000000000001100000000000000010000010010011",
72 => "0000000000000001000000000000001100000000000000010000010010101",
73 => "0000000000000001000000000000001100000000000000110000010010111",
74 => "0000000000000011000000000000100100000000000000110000010011001",
75 => "0000000000000001000000000000000100000000000000110000010011011",
76 => "0000000000000011000000000001001100000000000000110000010011110",
77 => "0000000000000001000000000000000100000000000000110000010100001",
78 => "0000000000000101000000000000001100000000001000110000010100011",
79 => "0000000000000001000000000000001100000000000000110000010100101",
80 => "0000000000000001000000000000001100000000001001000000010100111",
81 => "0000000000000001000000000000000100000000000000110000010101001",
82 => "0000000000000001000000000000100100000000000000110000010101011",
83 => "0000000000000001000000000000001100000000000000010000010101101",
84 => "0000000000101001000000000000001100000100010101000000010101111",
85 => "0000000000000001000000000000001100000000000000110000010110001",
86 => "0000000000000101000000000000001100000000000000110000010110011",
87 => "0000000000000001000000000000001100000000000000010000010110101",
88 => "0000000000001011000000000000001100000000010100010000010110111",
89 => "0000000010010011000000000000001100000000000000010000010111001",
90 => "0000000100100000000000000000010100000000000000110000010111011",
91 => "0000000000000001000000000000010100000000000000110000010111101",
92 => "0000000000000001000000000000001100000010001010000000010111111",
93 => "0000010001010101000000000100100100000000000000110000011000001",
94 => "0000000000000001000000000000000100000000000000110000011000011",
95 => "0000000000000001000000001000100100000000000000110000011000101",
96 => "0000000000000001000000000000001100000000000001010000011000111",
97 => "0000000000000001000000000000000100000000000000110000011001001",
98 => "0000000000000001000000000000001100000000000010010000011001011",
99 => "0000000000000001000000000000001100000000000010110000011001101",
100 => "0000000000000001000000000000001100000000000001010000011001111",
101 => "0000000000000001000000000000001100000000000000110000011010001",
102 => "0000000000000101000000000000001100000000000101010000011010011",
103 => "0000000000000001000000000000001100000000000001010000011010101",
104 => "0000001010000101000000000000001100000000000000010000011010111",
105 => "0000000000000001000000000000001100000000000001010000011011001",
106 => "0000000000000001000000000000000100000000000000110000011011100",
107 => "0000000001010001000000000000000100000000000000110000011011110",
108 => "0000000000001001000000000000000100000000000000110000011100000",
109 => "0000000000000001000000000000001100000000000010010000011100010",
110 => "0000000000000001000000000000001100000000000001010000011100101",
111 => "0000000000000001000000000000001100000000000000010000011101000",
112 => "0000000000000001000000000000001100000000010001000000011101010",
113 => "0000001000100000000000000000001100000000000000010000011101100",
114 => "0000000000000001000000000000001100000000000000010000011101110",
115 => "0000000000000001000000000000001100000000000000010000011110000",
116 => "0000001000101010000000000000001100000000000100010000011110010",
117 => "0000000000000001000000000000001100000000000000010000011110100",
118 => "0000000000101011000000000001000000000000000000110000011110110",
119 => "0010000100000001000000000000001100000000000000010000011111001",
120 => "0000000000000001000000000000001100000000000000010000011111011",
121 => "0000000000000001000000000000001100000000000000110000011111110",
122 => "0000000000000001000000000001000100000000000000110000100000001",
123 => "0000000000000001000000000000000100000000000000110000100000100",
124 => "0000000000000001000000000000000100000000000000110000100000110",
125 => "0000000000000001000000000000001100000001000000100000100001000",
126 => "0000000000000001000000000000000100000000000000110000100001010",
127 => "0000000000000001000000000000001100000000000000010000100001100",
128 => "0000000000000001000000000001000100000000000000110000100001110",
129 => "0000000000000001000000000000001100000000000001010000100010000",
130 => "0000000000000001000000000000001100000000000100010000100010010",
131 => "0000000000010011000000000000001100000000000000010000100010100",
132 => "0000000000001001000000000000001100000000100001010000100010110",
133 => "0000000000000001000000000000001100000000000000110000100011000",
134 => "0000000000000001000000000000000100000000000000110000100011010",
135 => "0000000000000001000000000000000100000000000000110000100011100",
136 => "0000000000000011000000000000001100000000010000110000100011110",
137 => "0000000000000001000000000000001100000000000010010000100100000",
138 => "0000001000001010000000000000001100000000001010010000100100010",
139 => "0000000001001010000000000000001100000010001000000000100100100",
140 => "0000000100000101000000000000001100000000000000110000100100110",
141 => "0000000000000011000000000000001100000000000000110000100101000",
142 => "0000000000000001000000101001000000000000000000110000100101010",
143 => "0000000000001011000000000000001100000000000000010000100101100",
144 => "0000000000000001000000000000001100000100100100100000100101110",
145 => "0000000000000001000000000000100100000000000000110000100110000",
146 => "0000000000000001000000000000000100000000000000110000100110010",
147 => "0000000000000001000000000000001100000000010000110000100110100",
148 => "0000000000000001000000000000001100000000000000010000100110110",
149 => "0000010101000001000000000000010100000000000000110000100111000",
150 => "0000000000000001000000010000100000000000000000110000100111010",
151 => "0000000000000001000000000000001100000000000000010000100111100",
152 => "0000000000000001000000000000000100000000000000110000100111110",
153 => "0000000000000101000000000000001100000000000001010000101000001",
154 => "0000000000000001000000000000001100000000000000010000101000011",
155 => "0000000000000001000000010000001000000000000000110000101000101",
156 => "0000000000000001000000000000001100000000000000010000101000111",
157 => "0000000000000001000000000000010100000000000000110000101001001",
158 => "0000000000000011000000000000001100000000000000010000101001011",
159 => "0000000000000001000000000000001100000000000000110000101001101",
160 => "0000000000000001000000000000000100000000000000110000101001111",
161 => "0000000000000001000000000000001100000000000000010000101010010",
162 => "0000000000000001000000000010000100000000000000110000101010100",
163 => "0000000000000101000000000000000100000000000000110000101010110",
164 => "0000000000000001000000000000001100000000000000010000101011000",
165 => "0000000000000001000000000000001100000000000100010000101011011",
166 => "0000000000000001000000000000001100000000000001010000101011101",
167 => "0000000000000001000000000000001100000000000000010000101011111",
168 => "0000000000000001000000010010100000000000000000110000101100001",
169 => "0000000010101011000000000000001100000000001010010000101100011",
170 => "0000000000000001000000000000001100000000001000010000101100101",
171 => "0000000000000101000000000000000100000000000000110000101100111",
172 => "0000000000000001000000000000001100000000001001000000101101001",
173 => "0000000000000011000000000000000100000000000000110000101101011",
174 => "0000000000000001000000000001010100000000000000110000101101101",
175 => "0000000000001001000000000000001100000000000000010000101101111",
176 => "0000000000000001000000000000001100000000000000110000101110001",
177 => "0000001000100101000000000010010100000000000000110000101110100",
178 => "0000000000000001000000000000001100000000000000010000101110111",
179 => "0000000000000001000000000000001100000000000000010000101111001",
180 => "0000000000001011000000000000010100000000000000110000101111011",
181 => "0000000000100011000000001001001000000000000000110000101111101",
182 => "0000000000000001000000000000001100000000010000100000101111111",
183 => "0000000000001011000000000000000100000000101000110000110000001",
184 => "0000000000000001000000000000001100000010010000000000110000011",
185 => "0000000000000001000000000000000100000000000000110000110000101",
186 => "0000000000000001000000000000001100000000000000010000110000111",
187 => "0000000000000001000000000000001100000000000000010000110001001",
188 => "0000000000010001000000000000001100000000000010110000110001100",
189 => "0000000100000001000000000000001100000000000000010000110001110",
190 => "0000001000001011000000000000001100000000000000010000110010000",
191 => "0000000000000001000000000000001100000000000000010000110010010",
192 => "0000000000000001000000010000101000000000000000110000110010100",
193 => "0000000000000001000000000000001100000000000001010000110010110",
194 => "0000000000000001000000000000001100000000000001010000110011000",
195 => "0000000000000001000000000000001100000000000000010000110011010",
196 => "0000000000000001000000000000000100000000000000110000110011100",
197 => "0000000000000001000000000000001100000000000000110000110011110",
198 => "0000000000000001000000100100010100000000000000110000110100000",
199 => "0000000000000001000000000001010100000000000000110000110100010",
200 => "0000000000010001000000000000001100000000000000010000110100100",
201 => "0000000100100010000000000000001100000000000100110000110100110",
202 => "0000000000000011000000000000001100000000000000110000110101000",
203 => "0000000000000001000000000000001100000000100100010000110101011",
204 => "0000000000000011000000000001001100000000000000110000110101101",
205 => "0000000000000001000000000000001100000000000000110000110101111",
206 => "0000010000010001000000000000010100000000000000110000110110001",
207 => "0000000000000001000000000000100100000000000000110000110110100",
208 => "0000000000000001000000000000001100000000001000010000110110111",
209 => "0000000000010001000000000000001100000000000000110000110111001",
210 => "0000000000000001000000000000100100000000000000110000110111011",
211 => "0000000000000001000000000000001100000000000000110000110111101",
212 => "0000000000000001000000000000001100000000000000110000110111111",
213 => "0000000000000011000000000000001100000000000000010000111000001",
214 => "0000000000000001000000000000001100000000101010100000111000011",
215 => "0000000000000001000000000000001100000000000000110000111000101",
216 => "0000010001010010000000000000001100000000000000110000111001000",
217 => "0000000000000001000000000000001100000000001001000000111001010",
218 => "0000000000000001000000000000001100000000000000010000111001101",
219 => "0000000000000001000000000000001100000000000000010000111001111",
220 => "0000000000000001000000100100001000000000000000110000111010001",
221 => "0000000000000001000000000000000100000000000000110000111010011",
222 => "0000000000000001000000000000001100000000000000010000111010101",
223 => "0000001000101000000000000000001100000000010000010000111010111",
224 => "0000000000000001000000000000001100000000000000010000111011010",
225 => "0000000000000001000000101000010100000000000000110000111011101",
226 => "0000000000000001000000000001001100000000000000110000111011111",
227 => "0000000000000011000000000000001100000010000101010000111100001",
228 => "0000000000000001000000010010101000000000000000110000111100011",
229 => "0000000000000011000000000000001100000000000000010000111100101",
230 => "0000000000000001000000000000000100000000000000110000111100111",
231 => "0000000000000001000000000000000100000000000000110000111101010",
232 => "0000000000000001000000000000000100000000000000110000111101100",
233 => "0000000000000011000000000000010100000000000000110000111101110",
234 => "0000000000000001000000000000001100000000000000010000111110000",
235 => "0000001000001000000000000000001100000000000000010000111110011",
236 => "0000000000000001000000000000001100000000000000110000111110110",
237 => "0000000000000001000000000000001100000000000100110000111111000",
238 => "0000000100000101000000000000000100000000000000110000111111010",
239 => "0000000000000001000000000000001100000000000000010000111111100",
240 => "0000000000000001000000000000000100000000000000110000111111110",
241 => "0000000000000001000000000000001100000000000000010001000000000",
242 => "0000000000000001000000000000001100000000000000010001000000011",
243 => "0001000100010010000000000000001100000000000001010001000000110",
244 => "0000000000000001000000000000000100000000000000110001000001000",
245 => "0000000000000001000000000100001100000000000000110001000001010",
246 => "0000000000000001000000000000100100000000000000110001000001100",
247 => "0000000000000001000000000000001100000000000000110001000001110",
248 => "0000000000000001000000000000000100000000000000110001000010000",
249 => "0000000000000001000000000000001100000000000100010001000010011",
250 => "0000000000000001000000000000000100000000000000110001000010110",
251 => "0000000000000011000000000000001100000000000000010001000011000",
252 => "0000000000000001000000000000001100000000000100110001000011010",
253 => "0000000000000001000000000000001100000001001010010001000011100",
254 => "0000000000000001000000000000001100000000000000010001000011110",
255 => "0000000000000001000000000000001100000010000001000001000100000",
256 => "0000000000000001000000000000100100000000000000110001000100011",
257 => "0000000000101011000000000000001100000000000000110001000100101",
258 => "0000000000000001000000000000001100000001000100010001000100111",
259 => "0000000000000001000000000000000100000000000000110001000101001",
260 => "0000001000100100000000000000001100000000100001010001000101011",
261 => "0000000000000001000000000101000100000000000000110001000101101",
262 => "0000000000000001000000000000001100000000000010110001000110000",
263 => "0000000000000000000000001010010100000000000000110001000110010",
264 => "0000000000000001000000000000001100000000000000010001000110100",
265 => "0000000000000001000000000000000100000000000000110001000110110",
266 => "0000000000001001000000000000001100000000000000010001000111000",
267 => "0000001010000011000000000000101100000000000000110001000111010",
268 => "0000000000000001000000001001000000000000000000110001000111100",
269 => "0000000000001001000000000000001100000000000000010001000111110",
270 => "0000000000000001000000000000001100000000000000010001001000000",
271 => "0000000000000001000000000000101100000000000000110001001000010",
272 => "0000000000000001000000000000001100000000000000010001001000100",
273 => "0000000000000001000000000000001100000000000000110001001000110",
274 => "0000000000000001000000000000000100000000000000110001001001000",
275 => "0000000000101001000000000001000100000000000000110001001001010",
276 => "0000000000000001000000000000001100000000000000110001001001100",
277 => "0000000000000001000000000000001100000000000000110001001001110",
278 => "0000000000000001000000001001010100000000000000110001001010000",
279 => "0000000000000001000000000000001100000000000000010001001010010",
280 => "0000000000001011000000000000010100000000000000110001001010100",
281 => "0000000000000001000000000000001100000000000000010001001010110",
282 => "0000000010010101000000000000001100000000000000110001001011000",
283 => "0000000000000011000000000000100100000000000000110001001011010",
284 => "0000000000000001000000000000001100000000000000010001001011100",
285 => "0000000000000001000000000000000100000000000000110001001011110",
286 => "0000000000000001000000000000000100000000000000110001001100000",
287 => "0000000000000001000000000000001100000000000000110001001100010",
288 => "0000000000000001000000000000001100000000000000010001001100100",
289 => "0000000000000001000000000000001100000000000000010001001100111",
290 => "0000000000000001000000000000001100000000000000010001001101001",
291 => "0000000000000001000000000000001100000000000100010001001101011",
292 => "0000000000000001000000000000001100000000000000110001001101110",
293 => "0000000000000001000000000000001100000000000000010001001110000",
294 => "0000000000000001000000000000000100000000000000010001001110010",
295 => "0000000000000001000000000000000100000000000000110001001110100",
296 => "0000000000000001000000000000001100000000101001000001001110110",
297 => "0000000000000001000000000000001100000000001010100001001111000",
298 => "0000000001010010000000000000001100000000101001010001001111010",
299 => "0000000000000001000000000000000100000000000000110001001111100",
300 => "0000000000000001000000000000001100000000000001010001001111110",
301 => "0000000000000001000000000000001100000000001010010001010000000",
302 => "0000000000000001000000000000001100000000000001010001010000010",
303 => "0000000000000001000000000000000100000000000000110001010000100",
304 => "0000000000000001000000000000001100000000000000110001010000110",
305 => "0000000000000001000000000000001100000000000000100001010001000",
306 => "0000000000000001000000000000001100000000000001010001010001010",
307 => "0000000000000001000000000000000100000000000000110001010001100",
308 => "0000000000000001000000000000001100000000000001010001010001110",
309 => "0000000000000101000000000000001100000000000000010001010010000",
310 => "0000000000000001000000000000001100000000000101010001010010010",
311 => "0000000000000001000000000000001100000000000001010001010010100",
312 => "0000000000000001000000000000101100000000000000110001010010110",
313 => "0000000000000001000000000000000100000000000000110001010011000",
314 => "0000000000000001000000000000000100000000000000110001010011010",
315 => "0000000000000001000000000000001100000000000000110001010011100",
316 => "0000000000000001000000000000001100000000101010000001010011110",
317 => "0000000000000001000000000000001100000000000000100001010100000",
318 => "0000000000000001000000000000000100000000000000110001010100011",
319 => "0001001010010101000000000000000100000000000000110001010100110",
320 => "0000000000000001000000001010000000000000000000110001010101001",
321 => "0000000000000001000000000000001100000000000101010001010101011",
322 => "0000000000000001000000000000001100000000000001010001010101101",
323 => "0001000010000010000000000000001100000000000010010001010101111",
324 => "0000000000000001000000000100000100000000000000110001010110001",
325 => "0000000000000001000000000000001100000000000000010001010110011",
326 => "0000000000010001000000000000001100000000100100110001010110101",
327 => "0000000000000001000000000000001100000000000000010001010110111",
328 => "0000000000000001000000000000010100000000000000110001010111010",
329 => "0000000000000001000000000000001100000000000000010001010111100",
330 => "0000000001001001000000000000000100000000000000110001010111110",
331 => "0000000000000001000000000000001100000000000000010001011000000",
332 => "0000000010010101000000000001010100000000000000110001011000010",
333 => "0000000000000001000000000000001100000000000010110001011000100",
334 => "0000000000000011000000000000001100000000000000010001011000110",
335 => "0000000000000001000000000000000100000000000000110001011001000",
336 => "0000000000010101000000000000001100000000000000010001011001010",
337 => "0000000000000001000000000000000100000000000000110001011001101",
338 => "0000000000000001000000000000001100000000000000110001011010000",
339 => "0000000001010010000000000000001100000000000000010001011010010",
340 => "0000000000000001000000000010100100000000000000110001011010100",
341 => "0000000000001001000000000000100100000000000000110001011010110",
342 => "0000000000100101000000000000001100000000000000010001011011000",
343 => "0000000000000011000000000000001100000000000000010001011011010",
344 => "0000010010000000000000000000000100000000000000110001011011100",
345 => "0000000000000001000000000000001100000000000000110001011011110",
346 => "0000000000000001000000000000001100000000001000110001011100000",
347 => "0000000000000001000000000000001100000000000000110001011100010",
348 => "0000001010101000000000000000000100000000000000110001011100100",
349 => "0000000000000001000000000000001100000000000000010001011100110",
350 => "0000000000000101000000000000001100000000000000010001011101000",
351 => "0000000000000011000000000100000000000000000000110001011101010",
352 => "0000000000000001000000000000001100000000000001010001011101100",
353 => "0000000000101011000000001000100100000000000000110001011101110",
354 => "0000000000000001000000000000000100000000000000110001011110000",
355 => "0000000000000001000000000000001100000000000100110001011110010",
356 => "0000000000000001000000000000101100000000000000110001011110100",
357 => "0000000000101001000000000000001100000000000100010001011110110",
358 => "0000000000000001000000000000001100000000100101010001011111000",
359 => "0000000000010011000000000000001100000000000000110001011111010",
360 => "0000000100100001000000000000001100000000000001010001011111101",
361 => "0000000000000001000000000000001100000000000000010001100000000",
362 => "0000000000000001000000000000001100000000000000110001100000011",
363 => "0000000000000101000000000000001100000000000000110001100000110",
364 => "0000000001001010000000000000001100000000101010110001100001001",
365 => "0000000000000001000000000000001100000000000001010001100001011",
366 => "0000000000000001000000000000000100000000000000010001100001101",
367 => "0000000000000001000000000000000100000000000000110001100010000",
368 => "0000000000000001000000000000001100000000000000010001100010011",
369 => "0000000000000001000000000000001100000000000000110001100010101",
370 => "0000000000000001000000000100100100000000000000110001100010111",
371 => "0000000000000001000000000000101100000000000000110001100011001",
372 => "0000000000000011000000000000000100000000000000110001100011011",
373 => "0000000000000001000000000000000100000000000000110001100011101",
374 => "0000010001000010000000000000001100000100000100010001100100000",
375 => "0000000000000001000000000000000100000000000000110001100100011",
376 => "0000000000000001000000000000001100000000000000010001100100110",
377 => "0000000000000001000000000000001100000000000000110001100101000",
378 => "0000000000000001000000000000000100000000000000110001100101010",
379 => "0000000000000001000000000000001100000000100010110001100101100",
380 => "0000000001001011000000000000001100000000000001010001100101110",
381 => "0000000000000001000000000000001100000000000000110001100110000",
382 => "0000000000000001000000000000001100000000000010110001100110010",
383 => "0000000000010101000000000000001100000010000100100001100110100",
384 => "0000000000000001000000000000001100000000000000010001100110110",
385 => "0000000001010011000000000000001100000000000000110001100111000",
386 => "0000000000000001000000000000001100000000000000110001100111010",
387 => "0000000000000001000000000000001100000000010010100001100111100",
388 => "0000000000000101000000001001000100000000000000110001100111110",
389 => "0000000000000101000000000000001100000100000100000001101000000",
390 => "0000000000000001000000000000001100000000000001010001101000010",
391 => "0000000000000001000000000000000100000000000000110001101000100",
392 => "0000000000000001000000000000000100000000000000110001101000110",
393 => "0000000010000011000000000000001100000000000000110001101001000",
394 => "0000000000000001000000000000001100000000000001010001101001010",
395 => "0000000000000001000000000000001100000000000000110001101001100",
396 => "0000000000000001000000000000001100000000000000010001101001110",
397 => "0000000001000101000000000000001100000000000000010001101010000",
398 => "0000000000010001000000000000001100000000000001010001101010010",
399 => "0000000000000001000000000000001100000000000000110001101010100",
400 => "0000000000000001000000000000010100000000000000110001101010110",
401 => "0000000000000001000000000000001100000000000000010001101011000",
402 => "0000000000000001000000000000000100000000000000110001101011010",
403 => "0000000000001001000000000000001100000000000000010001101011100",
404 => "0000000000000001000000000000001100000000000010010001101011110",
405 => "0000000000000001000000000000001100000000000000110001101100000",
406 => "0000000000001001000000000000001100000000000010010001101100010",
407 => "0000000000001001000000000000001100000000000100010001101100100",
408 => "0000000000000101000000000000001100000000000000010001101100110",
409 => "0000000000000001000000000000001100000000000000110001101101000",
410 => "0000000000000001000000000000001100000000000000110001101101010",
411 => "0000000000000001000000000000001100000000000000010001101101100",
412 => "0000000001001001000000000000001100000000000000110001101101110",
413 => "0000000000000001000000000000001100000000000000010001101110001",
414 => "0000000000000001000000000000000100000000000000110001101110011",
415 => "0000000000010011000000000001000100000000000000110001101110101",
416 => "0000000000001011000000000000010100000000000000110001101111000",
417 => "0000000000000001000000000000001100000000001000110001101111011",
418 => "0000000001010101000000000000001100000000000001010001101111101",
419 => "0000000000000001000000000000010100000000000000110001101111111",
420 => "0000000000001011000000000000001100000000000000110001110000001",
421 => "0000000000000001000000000000001100000000000000010001110000011",
422 => "0000000000000001000000000000001100000000000000010001110000101",
423 => "0000000100001000000000000000000100000000000000110001110000111",
424 => "0000000000000001000000000000000100000000000000110001110001001",
425 => "0000000000000001000000001000000100000000000000110001110001011",
426 => "0000000000000001000000000000001100000000000001010001110001101",
427 => "0000000000000001000000000000001100000000010000110001110001111",
428 => "0000000000000001000000000000000100000000000000110001110010001",
429 => "0000000000000001000000000100001100000000000000110001110010011",
430 => "0000000000000001000000000000001100000000000000010001110010101",
431 => "0000000000000001000000000101000100000000000000110001110010111",
432 => "0000000000000001000000000000001100000000000000110001110011001",
433 => "0000000000000001000000000000001100000000000000010001110011011",
434 => "0000000000000101000000000000010100000000000000110001110011101",
435 => "0000000000000001000000000000001100000000000000110001110011111",
436 => "0000000000000001000000000000000100000000000000110001110100001",
437 => "0000000000000001000000000000001100000000000000010001110100011",
438 => "0000000000000001000000000000001100000000000000110001110100101",
439 => "0000000010001011000000000000000100000000000000110001110100111",
440 => "0000000000000001000000000000001100000000000100000001110101001",
441 => "0000000000000001000000000000000100000000000000110001110101011",
442 => "0000000100000000000000000000001100000000000000010001110101101",
443 => "0000000000000001000000000000001100000000000000110001110101111",
444 => "0000000000000001000000000000000100000000000000110001110110001",
445 => "0000000000000001000000000000101000000000000001010001110110100",
446 => "0000000000001011000000000000001100000000000100110001110110110",
447 => "0000000000000111000000000000000100000000000000110001110111000",
448 => "0000000000000011000000000000001100000100010100100001110111010",
449 => "0000000000000001000000000000001100000000010010010001110111100",
450 => "0000000000000001000000000000001100000000000000110001110111110",
451 => "0000000000000001000000000000001100000000000000010001111000000",
452 => "0000000000000001000000000000000100000000000000110001111000011",
453 => "0000000000000011000000000000000100000000000000110001111000101",
454 => "0000000000000001000000000000001100000000000000010001111001000",
455 => "0000000000010011000000000000001100000000010010110001111001011",
456 => "0000000000000001000000000000000100000000000000110001111001101",
457 => "0000000000000001000000000000000100000000000001010001111001111",
458 => "0000000000000001000000000000001100000000000000010001111010001",
459 => "0000000000000001000000000000000100000000000000010001111010011",
460 => "0000000000000011000000000000001100000000000100110001111010110",
461 => "0000000000000001000000000000001100000000000100010001111011001",
462 => "0000000000000001000000000000001100000000000000110001111011100",
463 => "0000000000000001000000000000001100000000101000010001111011110",
464 => "0000000000000001000000000000001100000000000000110001111100001",
465 => "0000000000000001000000000000000100000000000000110001111100100",
466 => "0000000000000001000000000000001100000000000000110001111100110",
467 => "0000000000000001000000000000001100000000100100100001111101000",
468 => "0000000000000001000000001001001100000000000000110001111101010",
469 => "0000000000000001000000000000001100000000010000100001111101100",
470 => "0000000000000011000000000000001100000000000000010001111101110",
471 => "0000000000000001000000000000001100000000000000010001111110000",
472 => "0000000000000001000000000000001100000000000000110001111110010",
473 => "0000000000001001000000000000001100000000000000010001111110100",
474 => "0000000000000001000000001000010100000000000000110001111110111",
475 => "0000000000001001000000000000001100000000000000010001111111001",
476 => "0000000000000001000000000000000100000000000000110001111111011",
477 => "0000000000010101000000000000000100000000000000110001111111101",
478 => "0000000000000011000000000000001100000000100001010001111111111",
479 => "0000010000010100000000000000001100000000000000010010000000010",
480 => "0000000000000001000000000000000100000000000000110010000000100",
481 => "0000000000000001000000000000001100000000000100110010000000110",
482 => "0000000000000001000000000000000100000000000000110010000001001",
483 => "0000000000010011000000000001000000000000001000110010000001011",
484 => "0000000000000001000000100100001100000000000000110010000001101",
485 => "0000000000000001000000000000001100000000010100010010000001111",
486 => "0000000000000001000000000000001100000000000000110010000010001",
487 => "0000000000000001000000000000001100000000000000010010000010011",
488 => "0000000000000001000000000000001100000000000000110010000010101",
489 => "0000100001000100000000000001001100000000000000110010000010111",
490 => "0000000000000001000000000000001100000000000000010010000011001",
491 => "0000000000000001000000000000001100000000010000010010000011100",
492 => "0000000000000001000000000000001100000000000000010010000011110",
493 => "0000000000000001000000000000001100000000000000110010000100000",
494 => "0000001010000001000000000000001100000000000000010010000100010",
495 => "0000000000000001000000000000000100000000000000110010000100100",
496 => "0000000000000001000000000000001100000000000000110010000100110",
497 => "0000000000010101000000000000001100000000101001010010000101000",
498 => "0000000000000001000000000000001100000000001001010010000101010",
499 => "0000000000000001000000000000001100000010101000010010000101100",
500 => "0000000000000001000000000000001100000000010010110010000101110",
501 => "0000010100000100000000000000001100000000100010010010000110000",
502 => "0000000000000001000000000000000100000000000000110010000110010",
503 => "0000000000000001000000000000000100000000000000110010000110100",
504 => "0000000000000001000000000000001100000000000000010010000110110",
505 => "0000000000000001000000000000001100000000010001010010000111000",
506 => "0000100010010001000000000100101100000000000000110010000111010",
507 => "0000000000000001000000000000001100000000000000110010000111100",
508 => "0000000000000001000000000000001100000000000000110010000111110",
509 => "0000000000010011000000000001010100000000000000110010001000000",
510 => "0000000010010011000000001010000100000000000000110010001000010",
511 => "0000000000000001000000000000001100000000000000110010001000100",
512 => "0000000000000011000000000000001100000001000010010010001000110",
513 => "0000000000000001000000000000001100000000000100010010001001000",
514 => "0000000000000001000000000000000100000000000000110010001001010",
515 => "0000000000000001000000000000000100000000000000110010001001100",
516 => "0000000000000001000000000000001100000000000000010010001001110",
517 => "0000000000100001000000000000001100000000000000010010001010000",
518 => "0000010001010001000000000000101100000000000000110010001010010",
519 => "0000000000000001000000000000001100000000001001010010001010100",
520 => "0000000000000001000000010000100000000000000000110010001010110",
521 => "0000000000000001000000000000000100000000000000110010001011001",
522 => "0000000000010001000000000000001100000000000000010010001011100",
523 => "0000000000000001000001000100000000000000000000110010001011110",
524 => "0000000000001001000000000000001100000000000000010010001100000",
525 => "0000000000010001000000000000001100000000000000110010001100010",
526 => "0000000000000001000000000000000100000000000000010010001100101",
527 => "0000000000000001000000000000001100000000000000110010001100111",
528 => "0000000000000001000000000000001100000000000000110010001101001",
529 => "0000000000000001000000000000001100000000000000110010001101011",
530 => "0000001010000010000000000010001000000000000000010010001101110",
531 => "0000000000000001000000000000000100000000000000110010001110000",
532 => "0000010000101010000000000001010100000000000000110010001110010",
533 => "0000000000000001000000000000001100000000000000010010001110100",
534 => "0000000000000001000000000000000100000000000000110010001110110",
535 => "0000000000000001000000010000010000000000000000110010001111000",
536 => "0000000000000001000000000000001100000000000001010010001111010",
537 => "0000000000000001000000000000001100000000000000110010001111100",
538 => "0000000001010011000000000000000100000000000000110010001111110",
539 => "0000000000000001000000000000000100000000000000110010010000000",
540 => "0000000000000001000000000000001100000000000000010010010000010",
541 => "0000000000000001000000000000001100000000000000010010010000100",
542 => "0000000010000011000000000000000100000000000000110010010000110",
543 => "0000000000000101000000000000001100000000000000010010010001001",
544 => "0000000000000001000000000000000100000000000000110010010001011",
545 => "0000000000000001000000000000001100000000000000010010010001101",
546 => "0000000000000001000000000010000100000000000000110010010001111",
547 => "0000000000000001000000000000000100000000000000110010010010010",
548 => "0000000000000001000000000000001100000000000000010010010010100",
549 => "0000000000000001000000000000010100000000000000110010010010111",
550 => "0000000000000001000000000000001100000000001010010010010011010",
551 => "0000000000000001000000000101010100000000000000110010010011100",
552 => "0000000000000001000000000000001100000000000000010010010011110",
553 => "0000000000000001000000000000001100000000000101010010010100000",
554 => "0000000000000001000000000000000100000000000000110010010100010",
555 => "0000000000000001000000000000001100000000000000110010010100101",
556 => "0000000000000001000000000000101100000000000000110010010100111",
557 => "0000000000000001000000000000000100000000000000110010010101001",
558 => "0000000000000001000000000000001100000000001010110010010101011",
559 => "0000000000000001000000000000001100000000000001010010010101101",
560 => "0000000000000101000000000000001100000000001000010010010110000",
561 => "0000000000000101000000000000001100000000000000010010010110010",
562 => "0000000000000001000000000001001100000000000100100010010110100",
563 => "0000000000000001000000000000000100000000000000110010010110110",
564 => "0000000000000001000000000000000100000000000101010010010111000",
565 => "0000000000000001000000000000001100000000000010110010010111010",
566 => "0000000000000001000000000000001100000000000000010010010111100",
567 => "0000000001010101000000000000001100000000000000010010010111110",
568 => "0000000000000001000000000000001100000000000000110010011000000",
569 => "0000000000000001000000000000001100000000000000110010011000010",
570 => "0000000000000011000000000000001100000001000000100010011000100",
571 => "0000000000000001000000000000001100000000000000110010011000110",
572 => "0000000000000001000000000000001100000000001010110010011001000",
573 => "0000000000000001000000000000001100000000100001010010011001010",
574 => "0000000000100011000000000000000100000000000000110010011001100",
575 => "0000000000000001000000000000001100000000000000110010011001110",
576 => "0000000000000001000000000000001100000000000000010010011010000",
577 => "0001001000100001000000000100001000000000000000110010011010010",
578 => "0000000000000101000000000000000100000000000000110010011010100",
579 => "0000000000000001000000000000001100000000000000010010011010110",
580 => "0000000000000001000000000000001100000000000000110010011011000",
581 => "0000000000000001000000000000000100000000000000110010011011010",
582 => "0000000000000001000000000000001100000000000000010010011011100",
583 => "0000000000000001000000000000000100000000000000110010011011110",
584 => "0000000000000011000000000000001100000000000000010010011100000",
585 => "0000000000000001000000000000000100000000000000110010011100010",
586 => "0000000000000101000000000000001100000000000000010010011100100",
587 => "0000000000000011000000000000100000000000000000110010011100110",
588 => "0000000000000001000000000101001100000000000000110010011101001",
589 => "0000000000000001000000000000001100000000000000110010011101100",
590 => "0000000000000001000000000000001100000000000000110010011101110",
591 => "0000000000000001000000000000001100000000000000110010011110000",
592 => "0000000000000001000000000000001100000000000000010010011110011",
593 => "0000000000000001000000000000000100000000000000110010011110110",
594 => "0000000000000001000000000000001100000000000000110010011111000",
595 => "0000000000000001000000000000010100000000000000110010011111011",
596 => "0000000100000001000000000000001100000000001001010010011111110",
597 => "0000000000000011000000000000001100000100000010010010100000000",
598 => "0000000000000001000000000000001100000000100100010010100000010",
599 => "0000000000010001000000000000001100000000000001010010100000100",
600 => "0000000000000001000000000000000100000000000000110010100000110",
601 => "0000000000000001000000000000001100000000010101010010100001000",
602 => "0000000000000011000000000000001100000000000100010010100001010",
603 => "0000000000000001000000000001001100000000000000110010100001100",
604 => "0000000000000001000000000000001100000000000000010010100001110",
605 => "0000000000000001000000000000001100000000000000010010100010000",
606 => "0000000000000001000000000000000100000000000000110010100010010",
607 => "0000000000000001000000010001000100000000000000110010100010100",
608 => "0000000000000001000000000000001100000000000000110010100010110",
609 => "0000000000000001000000000000001100000000000001010010100011000",
610 => "0000000000000001000000000010010100000000000000110010100011010",
611 => "0000000000000001000000000001010100000000000000110010100011100",
612 => "0000000000000001000000000000001100000000000000110010100011110",
613 => "0000000000000001000000000000001100000000000000110010100100000",
614 => "0000000000000001000000000000000100000000000000110010100100010",
615 => "0000000000000001000000000000001100000000000000010010100100100",
616 => "0000000000000001000000000000001100000000000100010010100100110",
617 => "0000000000000001000000000000001100000000000000010010100101000",
618 => "0000000000000001000000000000001100000000000000010010100101010",
619 => "0000000000000001000000000000001100000000000000110010100101100",
620 => "0000000000000001000000000000000100000000000000110010100101110",
621 => "0000000000000001000000000000001100000000000000110010100110000",
622 => "0000000000000001000000000000001100000000000000010010100110010",
623 => "0000000000000001000000000000001100000000000100010010100110100",
624 => "0000000000001011000000000000001100000000000010010010100110110",
625 => "0000000001010011000000000100010100000000000000110010100111001",
626 => "0000000000000001000000000000001100000000000000110010100111100",
627 => "0000000000000001000000000000001100000000100001010010100111110",
628 => "0000000000000001000000000000001100000000100101010010101000000",
629 => "0000000000000001000000000000001100000000000000010010101000010",
630 => "0000000010010001000000000000001100000000000000010010101000100",
631 => "0000000000000001000000000000000100000000000000010010101000110",
632 => "0000000000000001000000000000000100000000000000110010101001000",
633 => "0000000000000001000000000000000100000000000000110010101001010",
634 => "0000000000000001000000000000001100000000000010010010101001100",
635 => "0000000000000001000000000000001100000000000000110010101001110",
636 => "0000000000000001000000000000001100000000000000110010101010000",
637 => "0000000000000001000000000000001100000000000000110010101010010",
638 => "0000000000000001000000000000001100000000000010010010101010100",
639 => "0000000000000001000000000000001100000000000000010010101010110",
640 => "0000000000000001000000000000001000000000000000110010101011000",
641 => "0000000000000001000000000000001100000000001010110010101011010",
642 => "0000000000000001000000000000001100000000000000110010101011100",
643 => "0000000000000001000000000000001100000000000000110010101011110",
644 => "0000000000000001000000000000001100000000000001010010101100000",
645 => "0000000000000001000000000000001100000000001000110010101100010",
646 => "0000000000000001000000000000001100000000000000110010101100100",
647 => "0000000000000001000000000000000100000000000100000010101100110",
648 => "0000010010000000000000000000001100000010001000000010101101000",
649 => "0000000000000001000000000000001100000000000101010010101101010",
650 => "0000000000000001000000000000000100000000000000110010101101100",
651 => "0000000010000001000000000000010100000000000000110010101101110",
652 => "0000000000000001000000000000001100000000000000110010101110000",
653 => "0000000000000001000000000000001100000000000000010010101110010",
654 => "0000000000001011000000000000001100000000000000110010101110100",
655 => "0000000000000001000000000000001100000000001001010010101110110",
656 => "0000000000000011000000000000001100000010001010010010101111001",
657 => "0000010100101010000000000000001100000000100100010010101111011",
658 => "0000000000000101000000000000010100000000000000110010101111101",
659 => "0000000000000001000000000000010100000000000000110010101111111",
660 => "0000000000000001000000000000001100000000000000110010110000010",
661 => "0000000000000001000000101000010000000000001000000010110000100",
662 => "0000000000001001000000000000001100000000000001010010110000110",
663 => "0000000000000011000000000000000100000000000000110010110001000",
664 => "0000000000000001000000000000000100000000000000110010110001010",
665 => "0000000000101001000000000000001100000000000100010010110001100",
666 => "0000000000000001000000000000001100000000000000110010110001111",
667 => "0000000000000001000000000000001100000000000000110010110010010",
668 => "0000000000000001000000000001001100000000000000110010110010100",
669 => "0000000000000001000000000000100100000000000000110010110010110",
670 => "0000000000000011000000000000001100000000000010010010110011000",
671 => "0000000000000001000000000000001100000000000000010010110011010",
672 => "0000000000001001000000000100000000000000000000110010110011100",
673 => "0000000000000001000000000000101100000000010000000010110011110",
674 => "0000000000000001000000000000000100000000000000110010110100000",
675 => "0000000000000001000000000000010100000000000000110010110100010",
676 => "0000000000001001000000000000001100000000000000110010110100101",
677 => "0000000000000001000000000000001100000000000000010010110100111",
678 => "0000000000000001000000000000001100000000000000110010110101001",
679 => "0000000000010101000000000000001100000000000000010010110101100",
680 => "0000000000000001000000000000010100000000000000110010110101111",
681 => "0000000000000001000000000000001100000000000000110010110110010",
682 => "0000000000000001000000000000001100000000000000110010110110100",
683 => "0000000000101001000000000000001100000000010001010010110110110",
684 => "0000000100001001000000000000010100000000000000110010110111001",
685 => "0000000000000001000000000000001100000000101010110010110111011",
686 => "0000000000000001000000000000001100000000000000110010110111101",
687 => "0000000000000001000000000000000100000000000100100010111000000",
688 => "0000000000000001000000000000001100000000000000110010111000010",
689 => "0000000000000001000000000000000100000000000000110010111000100",
690 => "0000000000001001000000000000001100000000000000010010111000110",
691 => "0000000000000001000000000000000100000000001000110010111001000",
692 => "0000000000000001000000000000000100000000000000110010111001011",
693 => "0000000000000001000000000000010100000000000000110010111001101",
694 => "0000000000000011000000000000001100000000000001010010111001111",
695 => "0000000100100001000000000000001100000000000000010010111010010",
696 => "0000000000010101000000000000001100000000000000110010111010100",
697 => "0000000000000001000000000000001100000010001010100010111010110",
698 => "0000000000000001000000000000100100000000000000110010111011000",
699 => "0000000010100101000000001000000100000000000000110010111011010",
700 => "0000000010010001000000000001010100000000000000110010111011101",
701 => "0000000000010001000000000000000100000000000000110010111100000",
702 => "0000000000000001000000000001001100000000000000110010111100010",
703 => "0000000000000011000000000000000100000000000000010010111100100",
704 => "0000000000000001000000000000001100000000000000010010111100110",
705 => "0000000100100011000000000000000100000000000100010010111101001",
706 => "0000000000000001000000000000000100000000000000110010111101100",
707 => "0000000000000001000000000000010100000000000000110010111101111",
708 => "0000000000010101000000000000000100000000000000110010111110001",
709 => "0000000000000001000000001010010000000000000000110010111110011",
710 => "0000000000010010000000000000001100000000010100100010111110101",
711 => "0000000000000001000000000000001100000000010010010010111110111",
712 => "0000000010000101000000000000001100000000000000010010111111001",
713 => "0000010001000100000000000000001100000000000010110010111111011",
714 => "0000000000000001000000000000001100000000000000010010111111101",
715 => "0000000000000001000000010101001000000000000000110010111111111",
716 => "0000000000000001000000000000001100000000000000010011000000001",
717 => "0000000000000001000000000000001100000000000000010011000000011",
718 => "0000000000001011000000000000001100000000000000110011000000101",
719 => "0000000000000001000000000000001100000000100000010011000000111",
720 => "0000000000000001000000000000001100000000001001010011000001001",
721 => "0000000010101011000000000000000100000000000000110011000001011",
722 => "0000000001010001000000000000001100000000000000010011000001101",
723 => "0000000000000001000000000000001100000000000000110011000010000",
724 => "0000000000000001000000000000001100000000000000010011000010010",
725 => "0000000000000001000000010010000000000000000000110011000010100",
726 => "0000000000010011000000000000010100000000000000110011000010110",
727 => "0000000000001011000000000000001100000000010000110011000011001",
728 => "0000000000000001000000000000101100000000000000010011000011011",
729 => "0000000000000001000000000000010100000000000000110011000011101",
730 => "0000000000000001000000000000001100000000100101000011000011111",
731 => "0000000000000001000000000000001100000000000001010011000100001",
732 => "0000000000000001000000000000000100000000000000110011000100011",
733 => "0000000000000001000000000000001100000000000010110011000100101",
734 => "0000000000000001000000000000001100000000000000010011000100111",
735 => "0000000000000001000000000000001100000000000000010011000101001",
736 => "0000000000000001000000000000000100000000000000110011000101011",
737 => "0000001001000000000000000001001100000000000000110011000101101",
738 => "0000000010101000000000000000001100000000000001010011000101111",
739 => "0000000000000001000000000000100100000000000000110011000110001",
740 => "0000000000000001000000000000001100000100001000000011000110011",
741 => "0000000000000001000000000000000100000000000000110011000110101",
742 => "0000000000000001000000000001000100000000000000110011000110111",
743 => "0000000000000001000000000000001100000000000000110011000111001",
744 => "0000000000000011000000000000101000000001000100110011000111011",
745 => "0000000000000001000000000000000100000000000000110011000111101",
746 => "0000000000000001000000001001001100000000000000110011000111111",
747 => "0000000000000001000000000000001100000000000000010011001000001",
748 => "0000000000000001000000000000000100000000000000110011001000011",
749 => "0000000000000001000000000000100100000000000000110011001000101",
750 => "0000000000000001000000000000001100000000000000110011001000111",
751 => "0000000000000011000000000000001100000000000000110011001001001",
752 => "0000000000000001000000000000001100000000101010100011001001100",
753 => "0000000000000001000000000000001100000000000000110011001001111",
754 => "0000000000000001000000000000001100000000000000010011001010001",
755 => "0000000000000001000000000000001100000000000000010011001010011",
756 => "0000000000000001000000100101000000000000000000110011001010101",
757 => "0000000000000001000000000000000100000000000000110011001011000",
758 => "0000000000000001000000000000001100000000000000110011001011011",
759 => "0000000000000001000000000000000100000000000000110011001011110",
760 => "0000000000000001000000000010101100000000000000110011001100000",
761 => "0000000000000001000000000000001100000000000000110011001100010",
762 => "0000000000000001000000000000001100000000101010010011001100101",
763 => "0000000000000011000000000000001100000001010100000011001100111",
764 => "0000000000001011000000000000010100000000000000110011001101001",
765 => "0000000000000001000000000000001100000000000000110011001101011",
766 => "0000000000000001000000000000001100000000000000010011001101101",
767 => "0000000000000001000000000000000100000000000000110011001101111",
768 => "0000000000000001000000001010100100000000000000110011001110001",
769 => "0000000000000001000000000000001100000000000000110011001110011",
770 => "0000000000000001000000000000001100000000000000010011001110101",
771 => "0000000000010001000000000000001100000000000000110011001111000",
772 => "0000000000000001000000000000001100000000000000110011001111010",
773 => "0000000000000001000000000000001100000000000010010011001111100",
774 => "0000000000000001000000000000101100000000000000110011001111110",
775 => "0000000000000001000000000000001100000000000000110011010000000",
776 => "0000000000000001000000000000101100000000000000000011010000011",
777 => "0000000000000001000000000000001100000000000000110011010000101",
778 => "0000000000000011000000001001010000000000000000110011010000111",
779 => "0000000000000001000000000000001100000000001000010011010001010",
780 => "0000000000000011000000000100001100000000000000110011010001100",
781 => "0000000000000001000000000000001100000000000000000011010001110",
782 => "0000000000000001000000000000001100000000000100110011010010000",
783 => "0000000000000001000000000000100100000000000000110011010010010",
784 => "0000000000000001000000010010010100000000000000110011010010100",
785 => "0000000000000101000000000000001100000000000000010011010010111",
786 => "0000010000100100000000000000001100000000000000110011010011001",
787 => "0000000000000001000000000001010100000000000000110011010011100",
788 => "0000000000000001000000000000000100000000000000110011010011110",
789 => "0000000000000001000000000000001100000000000000110011010100000",
790 => "0000000000000001000000000000000100000000000000110011010100010",
791 => "0000000000000101000000000000001100000000000000010011010100100",
792 => "0000000001000101000000000001000000000000000100110011010100110",
793 => "0000000000000001000000000000000100000000000000110011010101000",
794 => "0000000000000001000000000000001100000000000000010011010101010",
795 => "0000000000000001000000000000001100000000000000110011010101100",
796 => "0000000000000101000000000000010100000000100101010011010101110",
797 => "0000000000000001000000000000001100000000000000110011010110000",
798 => "0000000000000001000000000000001100000000000000010011010110010",
799 => "0000000000000001000000000000000100000000000000110011010110100",
800 => "0000000000000001000000000000001100000000000000110011010110110",
801 => "0000000000000001000000000000001100000000000000110011010111001",
802 => "0000000000000001000000000000001100000000000000110011010111011",
803 => "0000000000001001000000000000001100000000000000110011010111101",
804 => "0000000101010011000000000100000100000000000000010011010111111",
805 => "0000000000000001000000000000001100000000000000110011011000001",
806 => "0000000000000001000000000000010100000000000000110011011000011",
807 => "0000000000000001000000000000000100000000000000110011011000101",
808 => "0000000000000001000000000000001100000000000101010011011001000",
809 => "0000000000000001000000000000000100000000000000110011011001010",
810 => "0000000000000001000000000000001100000000000001010011011001100",
811 => "0000000000010011000000000000001100000000000010010011011001110",
812 => "0000000000000011000000000000001100000000000000010011011010000",
813 => "0000000000000001000000000010001100000000000000110011011010010",
814 => "0000000000000001000000000000001100000000001010010011011010100",
815 => "0000000000000001000000000001001100000000000000110011011010110",
816 => "0000000000000001000000000000000100000000000000010011011011000",
817 => "0000000000000001000000000000001100000000001000000011011011010",
818 => "0000000000000001000000010101001000000000000000110011011011100",
819 => "0000000000000001000000000000001100000000000000110011011011110",
820 => "0000000000100001000000000100000100000000000000010011011100001",
821 => "0000000000000001000000000000001100000000000000110011011100011",
822 => "0000000000000011000000000000001100000010001000000011011100101",
823 => "0000000000000001000000001000100100000000000000110011011100111",
824 => "0000000000000001000000000000000100000000000000110011011101001",
825 => "0000000000000001000000000000001100000000000000110011011101011",
826 => "0000000000001001000000000000001100000010010001000011011101101",
827 => "0000000000000001000000000000001100000000100000010011011101111",
828 => "0000000000000001000000000000001100000000000000010011011110001",
829 => "0000000000000011000000000000001100000000000000010011011110011",
830 => "0000000000000001000000000000001100000000000000010011011110101",
831 => "0000000000000001000000000000001100000000000000110011011110111",
832 => "0000000000000001000000000000001100000000000010110011011111001",
833 => "0000000000000001000000000000001100000000000000110011011111011",
834 => "0000000000000001000000000000000100000000000000010011011111110",
835 => "0000000000000001000000000000001100000000000000110011100000000",
836 => "0000000000000001000000000010001100000000000100100011100000010",
837 => "0000000000000001000000000000101100000000000000110011100000100",
838 => "0000000000000001000000000000001100000000100001010011100000110",
839 => "0000000000000001000000000000001100000000000000110011100001000",
840 => "0000000000000001000000000000001100000000000000110011100001010",
841 => "0000000000000001000000000000001100000000000000110011100001100",
842 => "0000000000000001000000000000001100000000000000010011100001110",
843 => "0000000000000001000000000000001100000000000100010011100010000",
844 => "0000000000000001000000000000001100000001000100000011100010010",
845 => "0000000000000101000000000000000100000000000000110011100010100",
846 => "0000000000000001000000000010101100000000000000110011100010110",
847 => "0000000000000001000000000000001100000000000000010011100011000",
848 => "0000000000000001000000000000000100000000000000110011100011010",
849 => "0000000000000001000000000000010100000000000000010011100011100",
850 => "0000000000000011000000000000001100000000000000110011100011110",
851 => "0000000000001001000000000000000100000000000000110011100100000",
852 => "0000000000000001000000000000001100000000000000010011100100011",
853 => "0000000000000001000000000000000100000000000000110011100100101",
854 => "0000000000000001000000000000001100000000000000110011100100111",
855 => "0000000000000001000000000000001100000000000000110011100101001",
856 => "0000000000000000000000000000010100000000000000110011100101100",
857 => "0000000000000011000000000000000100000000000000110011100101110",
858 => "0000000000000001000000000000001100000000000000110011100110000",
859 => "0000000000000001000000000000001100000000000000010011100110010",
860 => "0000000000000001000000000000010100000000000000110011100110101",
861 => "0000000000000001000000000010101100000000000000110011100110111",
862 => "0000000000000001000000000000001100000000000000110011100111010",
863 => "0000000000000001000000000000000100000000000000110011100111101",
864 => "0000000000000001000000000000010100000000000000110011100111111",
865 => "0000000000000001000000000000001100000000000000110011101000001",
866 => "0000000000000001000000000000001100000000000001010011101000100",
867 => "0000000000000011000000000000000100000000000000010011101000111",
868 => "0000010100010101000000000000001100000000000000010011101001001",
869 => "0000000000000001000000000000000100000000000000110011101001100",
870 => "0000000000000001000000000000101100000000000000110011101001110",
871 => "0000001010010001000000000000001100000000000001010011101010000",
872 => "0000000000000001000000000000001100000100000010010011101010010",
873 => "0000000000000001000000000000000100000000000000110011101010100",
874 => "0000000000000001000000000000001100000000000001000011101010110",
875 => "0000000000000001000000000100000100000000000100000011101011000",
876 => "0000000000000001000000000000000100000000000000110011101011010",
877 => "0000000100100010000000000000000100000000000000110011101011101",
878 => "0000000000000001000000000000001100000000000000110011101011111",
879 => "0000000000000001000000000000001100000000000000110011101100001",
880 => "0000000000000001000000000000001100000000000000110011101100011",
881 => "0000000010101011000000000000000100000000000000110011101100101",
882 => "0000000000001011000000000000001100000000000000110011101100111",
883 => "0000000000000001000000000000101100000000000000110011101101001",
884 => "0000000000000001000000000000001100000000000000110011101101011",
885 => "0000000000000001000000000000001100000000100101000011101101101",
886 => "0000000000000001000000000000100100000000000000110011101101111",
887 => "0000000000000001000000000000001100000000000000010011101110001",
888 => "0000000000000101000000000000001100000000000010010011101110011",
889 => "0000000000000001000000000000010100000000000001010011101110101",
890 => "0000000000000001000000000000000100000000000000110011101110111",
891 => "0000000000000001000000000001000100000000000000110011101111001",
892 => "0000000000000001000000000000000100000000000000110011101111011",
893 => "0000000000000101000000000000001100000000000000010011101111101",
894 => "0000010001000010000000000000001100000000000000110011101111111",
895 => "0000000000000001000000000000010100000000000000110011110000001",
896 => "0000000000000011000000000000001100000000100010000011110000011",
897 => "0000000000000001000000000000111100000000000000010011110000101",
898 => "0000000000001001000000000000001100000000000000010011110000111",
899 => "0000000000000011000000000000001100000000000000010011110001001",
900 => "0000000000000001000001001001010000000000000000110011110001011",
901 => "0000000000000001000000000000001100000000010010110011110001101",
902 => "0000000000000001000000000000010100000000000000110011110001111",
903 => "0000000000000001000000100100000100000000000000110011110010001",
904 => "0000000000010011000000000000001100000001001010110011110010011",
905 => "0000000000001101000000000101000100000000000000110011110010101",
906 => "0000000000000001000000000010101100000000000000110011110010111",
907 => "0000000000000001000000000000001100000000000000010011110011001",
908 => "0000000000000001000000000000001100000000001010000011110011011",
909 => "0000000000000011000000000000000100000000000000110011110011101",
910 => "0000000000000001000000000000001100000000000000010011110011111",
911 => "0000000000000001000000000000001100000000000000010011110100001",
912 => "0000000000100001000000000000001100000101000101000011110100100",
913 => "0000000000000001000000000000010100000000000000110011110100111",
914 => "0000000000000001000000000000001100000000000000110011110101001",
915 => "0000000000000001000000000000001100000000000000010011110101011",
916 => "0000000000000001000000000000000100000000000000110011110101101",
917 => "0000000000000001000000000000001100000000000000010011110101111",
918 => "0000000000000001000000000000001100000000000000110011110110001",
919 => "0000000010001010000000000000001100000000000000010011110110011",
920 => "0000000000000001000001000100010000000000000000110011110110101",
921 => "0000000000000001000000000000001100000000000000110011110111000",
922 => "0000000000000001000000000000001100000000001000110011110111010",
923 => "0000000000100001000000010000010000000000000000110011110111100",
924 => "0000000000000001000000000000001100000000000000110011110111110",
925 => "0000000000000001000000000000001100000000000010110011111000000",
926 => "0000000000000001000000000000001100000000000000110011111000010",
927 => "0000000000000001000000010101001000000000000000010011111000100",
928 => "0000000000000001000000000000001100000000000000010011111000110",
929 => "0000000000000001000000000000001100000000000001010011111001000",
930 => "0000000000000001000000000000001100000000000000110011111001010",
931 => "0000000000000001000000000000100100000000010000000011111001100",
932 => "0000000000000001000000000000001100000000000000110011111001110",
933 => "0000000000000001000000000000001100000000000001010011111010000",
934 => "0000000000000001000000000000001100000000000000010011111010010",
935 => "0000000000000001000000000000000100000000000000010011111010100",
936 => "0000000000000101000000000000001100000000000000110011111010110",
937 => "0000000000000001000000000000001100000000000000110011111011000",
938 => "0000000000000001000000000010000100000000000000110011111011010",
939 => "0000000000000001000000000000001100000001000001000011111011100",
940 => "0000000000000011000000000000001100000000000000110011111011110",
941 => "0000000000010001000000000000001100000000000000010011111100000",
942 => "0000000000000001000000000000001100000000001000100011111100010",
943 => "0000000000000001000000000000001100000000000000010011111100100",
944 => "0000000000000001000000000000010100000000000000110011111100110",
945 => "0000000000000001000000000000001100000000000000110011111101000",
946 => "0000000000000001000000000000000100000000000000110011111101010",
947 => "0000000000000011000000000000001100000000000000110011111101101",
948 => "0000000000000001000000000000001100000000001000010011111110000",
949 => "0000000000000001000000000001001100000000000000110011111110010",
950 => "0000000000000001000000000000001100000000000000010011111110101",
951 => "0000000000000001000000000000001100000001001001010011111111000",
952 => "0000000000000001000000000000001100000000000000110011111111011",
953 => "0000000000000001000000000000000100000000000000110011111111101",
954 => "0000000000000001000000000000001100000000000000110100000000000",
955 => "0000000000000011000000000000101100000000000000110100000000010",
956 => "0000000000000001000000000000001100000000000000110100000000101",
957 => "0000000000000001000000000000010100000000000000110100000000111",
958 => "0000000000000001000000000000001100000000000000010100000001010",
959 => "0000000000000001000000000000001100000000000001010100000001100",
960 => "0000000000000011000000000000001100000000000000110100000001111",
961 => "0000000000000001000000000000000100000000000000110100000010001",
962 => "0000010000101010000000000000001100000000000001010100000010011",
963 => "0000000001010000000000000000001100000000000000110100000010110",
964 => "0000000000000001000000000000001100000000010001010100000011000",
965 => "0000000000000001000000000000001100000000000100010100000011010",
966 => "0000000000000001000000000000000100000000000000110100000011101",
967 => "0000000000000101000000000000000100000000000001010100000100000",
968 => "0000000000000001000000000000001100000000000000110100000100010",
969 => "0000000000000001000000000000000100000000000000010100000100101",
970 => "0000000000000001000000000000001100000000000000110100000100111",
971 => "0000000000001011000000000000101100000000000000010100000101001",
972 => "0000000001010011000000000000001100000000000000010100000101011",
973 => "0000000000000001000000101010001000000000000000110100000101101",
974 => "0000000000000001000000000000001100000000000001010100000101111",
975 => "0000000000000001000000000000001100000010010010010100000110001",
976 => "0000000000001011000000000000001100000010010100100100000110011",
977 => "0000000100000010000000000000001100000000000000010100000110101",
978 => "0000000000000001000000100000100000000000000000110100000111000",
979 => "0000000000101001000000000000001100000000000010010100000111011",
980 => "0000000000000001000000000000000100000000000000010100000111101",
981 => "0000000000000001000000000000000100000000000000110100001000000",
982 => "0000000000000001000000000000001100000000000000010100001000011",
983 => "0000000000000001000000000000001100000000000000010100001000101",
984 => "0000000000000001000000000000001100000000000000110100001000111",
985 => "0000000000000001000000000100101100000000000000110100001001001",
986 => "0000000000000001000000000000001100000000000000110100001001011",
987 => "0000000000000001000000000000001100000000000001010100001001101",
988 => "0000000000000001000000000000001100000000000000010100001001111",
989 => "0000000010010011000000000000001100000000000000110100001010001",
990 => "0000000000000001000000000000001100000000000000010100001010011",
991 => "0000000000000001000000000000001100000000000000110100001010110",
992 => "0000000000000001000000000100010100000000000000110100001011001",
993 => "0000000001000011000000000100010000000000000000110100001011011",
994 => "0000000000000001000001001001000000000000001010010100001011101",
995 => "0000000000000001000000000000001100000000000100110100001011111",
996 => "0000000000100001000000000000001100000000000101010100001100001",
997 => "0000000000000001000000000001001100000000000000110100001100011",
998 => "0000001000000011000000000000010100000000000000110100001100101",
999 => "0000000000000001000000000000101100000000000000110100001100111",
1000 => "0000000000000011000000000000001100000000000100110100001101001",
1001 => "0000000000010001000000000000001100000000100000010100001101011",
1002 => "0000000000000001000000000000100100000000000000110100001101101",
1003 => "0000000000000101000000000000001100000000000000110100001101111",
1004 => "0000000000000011000000000000000100000000000000110100001110001",
1005 => "0000000000000001000000000000001100000000000000110100001110011",
1006 => "0000000000000001000000000000001100000000001010010100001110101",
1007 => "0000000101001010000000000000001100000000000000110100001110111",
1008 => "0000000000000001000000000000001100000000000000010100001111001",
1009 => "0000000000000011000000000000001100000000000000010100001111011",
1010 => "0000000000000001000000000000001100000000001001010100001111110",
1011 => "0000000000000001000000000101000100000000000000110100010000000",
1012 => "0000000000000001000000000101001100000000000000110100010000010",
1013 => "0000000000000011000000000000001100000010001010100100010000101",
1014 => "0000000000000010000000000000001100000000001010110100010001000",
1015 => "0000000000000001000000000000001100000000000000110100010001010",
1016 => "0000000000000001000000000000000100000000000000110100010001100",
1017 => "0000000000100101000000000000001100000000000000010100010001111",
1018 => "0000000000000001000000000000010100000000000000110100010010010",
1019 => "0000000000101011000000000000001100000000000000110100010010101",
1020 => "0000000000000001000000000000001100000000000000010100010010111",
1021 => "0000000000000001000000000000001100000000000000110100010011001",
1022 => "0000000000001011000000000000001100000000000000010100010011100",
1023 => "0000000000001001000000000000001100000000000000010100010011110",
1024 => "0000000000001011000000000000001100000000000000110100010100000",
1025 => "0000000000000101000000000000001100000000000000010100010100010",
1026 => "0000000000000101000000000000001100000001010101000100010100100",
1027 => "0000000000000001000000000000001100000000000000110100010100110",
1028 => "0000000000100000000000000000001100000000000000010100010101000",
1029 => "0000000000000001000000000000001100000000000000110100010101010",
1030 => "0000000000000001000000000000001100000000000010110100010101100",
1031 => "0000000000000011000000000000001100000000000000110100010101110",
1032 => "0000000000000001000000000000001100000000100001000100010110000",
1033 => "0000000000000001000000000000001100000000000000010100010110010",
1034 => "0000000000000001000000000000010100000000000000110100010110100",
1035 => "0000000000000001000000000000001100000000000000010100010110110",
1036 => "0000000000000011000000000000001100000000000010010100010111000",
1037 => "0000000000000001000000000000001100000000000100100100010111010",
1038 => "0000000000000001000000000000000100000000000000110100010111100",
1039 => "0000000000000001000000000000001100000000000001010100010111110",
1040 => "0000000000000001000000000111010100000000000000010100011000000",
1041 => "0000000000000001000000000000000100000000000000110100011000010",
1042 => "0000000000100101000000000000101000000000000000010100011000100",
1043 => "0000000000000001000000000000000100000000000000110100011000110",
1044 => "0000000000000001000000001010100000000000000000110100011001000",
1045 => "0000000000000001000000000000001100000000000000100100011001011",
1046 => "0000000000000001000000000000001100000000000000010100011001101",
1047 => "0000000000000001000000000000001100000000000000110100011010000",
1048 => "0000000000000001000000000000001100000000000000010100011010011",
1049 => "0000000000000001000000001010100100000000000000110100011010101",
1050 => "0000000000000001000000000000000100000010001000000100011010111",
1051 => "0000000000000001000000000000010100000000000000110100011011001",
1052 => "0000000000000001000000001000001100000000000000110100011011011",
1053 => "0000000000000001000000000000001100000000000000110100011011101",
1054 => "0000000000001001000000000000001100000000000000010100011011111",
1055 => "0000000000000001000000000000001100000000001010100100011100001",
1056 => "0000000000000001000000000000001100000010100010000100011100011",
1057 => "0000000000000001000000000000001100000000000010010100011100101",
1058 => "0000000000000001000000000100010100000000000000110100011101000",
1059 => "0000000000000001000000000000001100000000000010110100011101011",
1060 => "0000000001000101000000000000010100000000000000110100011101101",
1061 => "0000000000000101000000000000001100000000001000010100011101111",
1062 => "0000000000000001000000000000001100000000000010010100011110001",
1063 => "0000000000000011000000000000001100000000101000010100011110011",
1064 => "0000000000000101000000000000000100000000000000110100011110101",
1065 => "0000000000010001000000000000001100000000000000110100011110111",
1066 => "0000000000000001000000000000010100000000001000100100011111001",
1067 => "0000000000000011000000000000001100000000000000010100011111011",
1068 => "0000000000101011000000000000000100000000000000110100011111101",
1069 => "0000000000000001000000010000000000000000000000110100011111111",
1070 => "0000000000000001000000000000001100000000010000110100100000001",
1071 => "0000000000000001000000000000001100000000000000110100100000011",
1072 => "0000000000000001000000000000001100000000000000110100100000101",
1073 => "0000000100100011000000000000001100000000000100010100100000111",
1074 => "0000000000000001000000000000001100000000000010110100100001001",
1075 => "0000000000000001000000000000000100000000000000110100100001100",
1076 => "0000000000000001000000000000000100000000000000110100100001110",
1077 => "0000000000000001000000000000001100000000000000110100100010000",
1078 => "0000000000000001000000000000000100000000000000110100100010010",
1079 => "0000000000000011000000000000001100000000001000010100100010100",
1080 => "0000000000010101000000000000000100000000000000110100100010110",
1081 => "0000000000000001000000000000001100000000000000110100100011001",
1082 => "0000000000000001000000000000001100000000000000010100100011100",
1083 => "0000000000000001000000000000001100000000000000010100100011110",
1084 => "0000000000000001000000000000001100000000000000010100100100001",
1085 => "0000000000000101000000000000001100000000000000010100100100011",
1086 => "0000000000000001000000000000000100000000000000110100100100101",
1087 => "0000000000000001000000000000000100000000000000110100100100111",
1088 => "0000000000000001000000000000001100000000000000010100100101010",
1089 => "0000000000000101000000000000001100000000000000110100100101100",
1090 => "0000000000000001000000000000000100000000000011110100100101110",
1091 => "0000000000000001000000000010001100000000000000110100100110000",
1092 => "0000000000000101000000000000001100000000000010110100100110010",
1093 => "0000000000000011000000000000001100000000000001010100100110100",
1094 => "0000000000000001000000000010010100000000000000010100100110110",
1095 => "0000000000000101000000000000001100000000000000010100100111001",
1096 => "0000000000000001000000000000001100000000010100010100100111100",
1097 => "0000000000000001000000000000001100000000000000110100100111111",
1098 => "0000000000000001000000000000000100000000000000110100101000001",
1099 => "0000000000000001000000000000001100000000000001010100101000100",
1100 => "0000000000000001000000000000000100000000000000110100101000110",
1101 => "0000000000000001000000000000001100000000000000110100101001001",
1102 => "0000000000000001000000000000001100000000000000010100101001011",
1103 => "0000010010010010000000001001000100000000000000110100101001101",
1104 => "0000000000000001000000000000001100000000000000010100101001111",
1105 => "0000000000000001000000000000001100000000000000110100101010001",
1106 => "0000000000000001000000000000010100000000000100010100101010011",
1107 => "0000000000000001000000000000001100000000000000110100101010101",
1108 => "0000000000000001000000001010000000000000000000110100101010111",
1109 => "0000000000001001000000000000001100000000000100110100101011001",
1110 => "0000000000000001000000000000000100000000000000110100101011011",
1111 => "0000000101000010000000000000001100000000000000010100101011101",
1112 => "0000000000010101000000000000001100000000000010110100101011111",
1113 => "0000000000000001000000000000001100000000000000010100101100001",
1114 => "0000000000000001000000000000000100000000000000110100101100011",
1115 => "0000000000000001000000000000001100000000000000110100101100101",
1116 => "0000000000001011000000000000001100000000000000010100101100111",
1117 => "0000000000000001000000000000001100000000000000010100101101001",
1118 => "0000000000000001000000000000010100000000000000110100101101011",
1119 => "0000000000000001000000000000001100000000001001010100101101101",
1120 => "0000001010001001000000000000010100000000000000110100101101111",
1121 => "0000000000000001000000000010101000000000000000110100101110001",
1122 => "0000000000000001000000000000000100000000000000100100101110011",
1123 => "0000000000000001000000000000000100000000000000110100101110101",
1124 => "0000000000000001000000000000001100000000000000110100101110111",
1125 => "0000000000000001000000000000001100000000000001010100101111001",
1126 => "0000000000000001000000000000000100000000000000110100101111011",
1127 => "0000000000000001000000000000000100000000000000110100101111101",
1128 => "0000000000000001000000000000010100000000000000110100101111111",
1129 => "0000000000000001000000000000001100000000000000110100110000001",
1130 => "0000000000000011000000000000101100000000000000110100110000011",
1131 => "0000000000000001000000100000100000000000000000110100110000101",
1132 => "0000000000100001000000000000001100000000000100010100110000111",
1133 => "0000000000000001000000000000001100000000000010010100110001001",
1134 => "0000000000000001000000000001000100000000000000010100110001011",
1135 => "0000000000000011000000000000001100000000010000100100110001101",
1136 => "0000000000000001000000000000000100000000000000110100110001111",
1137 => "0000000000000001000000000000001100000000010000010100110010001",
1138 => "0000000000000001000000000000001100000000000010010100110010100",
1139 => "0000000000000001000000000000001100000000000000110100110010111",
1140 => "0000000000000001000000000000001100000000101000010100110011010",
1141 => "0000000000000001000000000000001100000000000000010100110011100",
1142 => "0000000000000001000000000000001100000000101000100100110011111",
1143 => "0000000101000101000000000000001100000000000000010100110100001",
1144 => "0000000000000001000000000000010100000000000000010100110100011",
1145 => "0000000000000001000000000000000100000000000000110100110100101",
1146 => "0000000000000001000000000000001100000000000100110100110100111",
1147 => "0000000000000001000000000000001100000000000000110100110101001",
1148 => "0000000000001011000000000000001100000000000000110100110101011",
1149 => "0000000000000001000000000000001100000000000000110100110101101",
1150 => "0000000000000001000000000000001100000000000100110100110101111",
1151 => "0000000000000001000000000000001100000000001001010100110110001",
1152 => "0000000000100101000000000000001100000000000000010100110110011",
1153 => "0000000000000001000000000010010100000000000000110100110110101",
1154 => "0000000000000001000000000000001100000000000000010100110110111",
1155 => "0000000000000001000000000000001100000000100010100100110111001",
1156 => "0000000000000001000000000000001100000000000000110100110111011",
1157 => "0000000000000001000000000000000100000000000000110100110111101",
1158 => "0000000000000001000000000000001100000000000000010100110111111",
1159 => "0000000000000001000000000000001100000000000000110100111000001",
1160 => "0000000000000101000000000000000100000000000000110100111000011",
1161 => "0000000000000001000000000000001100000000000000010100111000101",
1162 => "0000000000000001000000000000010100000000000100010100111001000",
1163 => "0000000000000001000000000000001100000001000101000100111001010",
1164 => "0000000000000001000000000000001100000000000000110100111001100",
1165 => "0000000000000001000000000000001100000000000010010100111001110",
1166 => "0000000000000001000000000000001100000000000000010100111010000",
1167 => "0000001000001000000000000000001100000000000010010100111010010",
1168 => "0000000000001001000000000000001100000000000000010100111010100",
1169 => "0000000000000001000000001000001100000000000000110100111010110",
1170 => "0000000000000001000000000000001100000000100100010100111011000",
1171 => "0000000000000001000000000000001100000000000000110100111011010",
1172 => "0000010010010101000000000000000100000000000000110100111011100",
1173 => "0000000000000001000000000000001100000000000000010100111011110",
1174 => "0000000000000001000000000000001100000000000000110100111100000",
1175 => "0000000000000001000000000000001100000000000000110100111100010",
1176 => "0000000000000001000000000000000100000000000000110100111100100",
1177 => "0000000000000001000000000000001100000000000000110100111100110",
1178 => "0000000000000001000000000000001100000000000000110100111101001",
1179 => "0000000000001011000000000000001100000000000000110100111101011",
1180 => "0000000101000101000000000000001100000000000001010100111101110",
1181 => "0000000000000001000000000000001100000000000000110100111110001",
1182 => "0000100000100010000000000000000100000000000000110100111110100",
1183 => "0000000000000011000000000000000100000000000000110100111110110",
1184 => "0000000000000001000000000000010100000000001000100100111111000",
1185 => "0000000000000001000000000000001100000000000000110100111111011",
1186 => "0000000000000001000000000001000100000000000000010100111111101",
1187 => "0000000001000011000000000000001100000000000010010100111111111",
1188 => "0000000000000001000000000000001100000000000000110101000000001",
1189 => "0000000000000001000000000000000100000000000000110101000000011",
1190 => "0000000000000001000000000000001100000000000000110101000000101",
1191 => "0000000000000001000000000000001100000000000000110101000000111",
1192 => "0000000000000001000000000000001100000001000010000101000001001",
1193 => "0000000000000001000000000000001100000001000010100101000001011",
1194 => "0000000000000001000000000000001100000000000100110101000001101",
1195 => "0000000000000001000000000000001100000000000000110101000001111",
1196 => "0000000000000001000000000000001100000000000001010101000010001",
1197 => "0000000000000011000000000000001100000000000000110101000010011",
1198 => "0000000000000001000000000000001100000000000001010101000010101",
1199 => "0000000000000001000000000000000100000000000000110101000010111",
1200 => "0000000000000001000000000000001100000000000000010101000011001",
1201 => "0000000000000001000000000000001100000000000010000101000011011",
1202 => "0000000000000001000000000000000100000000000000110101000011101",
1203 => "0000000000000001000000000000001100000000000000110101000011111",
1204 => "0000000000000001000000000000100100000000000000110101000100001",
1205 => "0000000000000001000000000000001100000000000000110101000100011",
1206 => "0000000000000001000000100101010100000000000000110101000100101",
1207 => "0000001000101001000000000000001100000000000000110101000100111",
1208 => "0000000000000101000000000000010100000000000000110101000101001",
1209 => "0000000000000001000000100001000000000000000000110101000101011",
1210 => "0000000000000001000000000000001100000000000000010101000101110",
1211 => "0000000000000001000000000000001100000000000000110101000110001",
1212 => "0000000000000001000000000000001100000000000000010101000110100",
1213 => "0000000000000001000000000100001100000000000000110101000110111",
1214 => "0000000000000001000000000001000100000000000000110101000111001",
1215 => "0000000000000011000000000000001100000000000000010101000111011",
1216 => "0000000000000011000000000000001100000000000000010101000111101",
1217 => "0000000000001001000000000000001100000000000000010101000111111",
1218 => "0000100100100100000000000101010000000001010000010101001000001",
1219 => "0000000010010011000000000000001100000000000000010101001000011",
1220 => "0000000000000001000000000000001100000000101000100101001000101",
1221 => "0000000000000001000000000000001100000000000000110101001000111",
1222 => "0000000000000011000000000000001100000000000000110101001001001",
1223 => "0000000000000001000000000000001100000000000000110101001001011",
1224 => "0000000000000001000000000000001100000000000010110101001001101",
1225 => "0000000000000001000000000000001100000000000000010101001001111",
1226 => "0000000000000001000000000000001100000000000000010101001010001",
1227 => "0000000000000011000000000000001100000000000000110101001010100",
1228 => "0000000000000001000000000001000100000000000000110101001010110",
1229 => "0000000000000001000000000000001100000000000101000101001011000",
1230 => "0000000000000001000000000000101100000000000000110101001011010",
1231 => "0000000000000001000000000000010100000000000000110101001011100",
1232 => "0000000000000001000000000001001100000000000000110101001011110",
1233 => "0000000000000001000000000000001100000000000000010101001100000",
1234 => "0000000000000011000000000000000100000000000000110101001100011",
1235 => "0000000000000001000000000000000100000000000000110101001100110",
1236 => "0000000000000001000000001000101000000000000000110101001101000",
1237 => "0000000000000001000000000000001100000000001000110101001101010",
1238 => "0000000000000001000000010100100000000000000000110101001101100",
1239 => "0000000000001011000000000000001100000001000100010101001101111",
1240 => "0000000000000011000000001010000000000000000000110101001110001",
1241 => "0000000000000001000000000000001100000000000101010101001110011",
1242 => "0000000001010101000000001010101000000000000000110101001110101",
1243 => "0000000010010001000000000000001100000001010001000101001110111",
1244 => "0000000000000011000000000000010100000000000000110101001111010",
1245 => "0000000000000001000000000100100100000000000000110101001111100",
1246 => "0000000000000001000000100100100000000000000000110101001111110",
1247 => "0000000000000001000000000000001100000000000000010101010000000",
1248 => "0000000000000001000000000000000100000000000000110101010000010",
1249 => "0000000000000001000000000000001100000000000000010101010000100",
1250 => "0000000001001011000000000000001100000000000000010101010000110",
1251 => "0000000001000001000000000000001100000000000001010101010001000",
1252 => "0000000000000001000000000000000100000000000000110101010001010",
1253 => "0000000000000001000000000000001100000000000010010101010001100",
1254 => "0000000000000001000000000001000000000000000000110101010001110",
1255 => "0000000000000001000000000000000100000000000000110101010010000",
1256 => "0000000000000001000000000000010100000000000000110101010010010",
1257 => "0000000000000001000000000000001100000000000000010101010010101",
1258 => "0000000000000001000000000000001100000000000001010101010010111",
1259 => "0000000000000001000000000000001100000000001010010101010011001",
1260 => "0000000000000001000000000000001100000000000100110101010011011",
1261 => "0000000000000011000000000000001100000001010100010101010011101",
1262 => "0000000000101001000000000000001100000000000000010101010011111",
1263 => "0000000000000001000000000000001100000000000000110101010100010",
1264 => "0000000000000001000000000000000100000000000000110101010100100",
1265 => "0000000000000001000000010010100100000000000000110101010100111",
1266 => "0000000000000111000000000000001100000000000000110101010101010",
1267 => "0000000000000001000000000000000100000000000000110101010101101",
1268 => "0000000000000001000000000000000100000000000000110101010101111",
1269 => "0000010001010010000000000100101100000000000000110101010110001",
1270 => "0000000000000001000000000000001100000000000001010101010110011",
1271 => "0000000000000001000000000000001100000000000000010101010110101",
1272 => "0000000000000001000000000000001100000000001010010101010110111",
1273 => "0000000000000001000000000000101100000000000000110101010111001",
1274 => "0000000000000001000000000000001100000000000000110101010111011",
1275 => "0000000000000011000000000000000100000000000000110101010111101",
1276 => "0000000000000101000000000000001100000000000000110101010111111",
1277 => "0000000000000001000000000000000100000000000000110101011000001",
1278 => "0000000000000101000000000000001100000000000001010101011000011",
1279 => "0000000000000001000000000000001100000000000100010101011000101",
1280 => "0000000000000001000000000000001100000000000000110101011000111",
1281 => "0000000000000001000000000000001100000000000000010101011001001",
1282 => "0000000000000001000000000000001100000000000101010101011001011",
1283 => "0000000000000001000000000000001100000000000000110101011001101",
1284 => "0000000000000001000000010100000100000000000000110101011001111",
1285 => "0000001000000010000000000000000100000000000000110101011010001",
1286 => "0000000000000001000000000000001100000000000000110101011010011",
1287 => "0000000000000001000000000000001100000000000001010101011010101",
1288 => "0000000101000000000000000010100000000000000000110101011010111",
1289 => "0000000000000001000000000000101100000000000000110101011011001",
1290 => "0000000000000001000000000000001100000000000000110101011011100",
1291 => "0000000000000001000000000000000100000000000010110101011011110",
1292 => "0000000101000000000000000000001100000000000001010101011100001",
1293 => "0000000000000001000000000000001100000000000010010101011100011",
1294 => "0000000000000011000000000000001100000000000010110101011100110",
1295 => "0000000000000001000000000000001100000000000000010101011101000",
1296 => "0000000000000001000000000000001100000000000000110101011101011",
1297 => "0000000000000001000000000000010100000000000000110101011101101",
1298 => "0000001000000100000000000000001100000000000000110101011110000",
1299 => "0000000000000001000000000000001100000000001001010101011110011",
1300 => "0000000000000001000000000000001100000000000001010101011110110",
1301 => "0000000000000011000000000000000100000000000000110101011111000",
1302 => "0000010101000100000000000000001100000001000000010101011111011",
1303 => "0000000000000001000000000000000100000000000000110101011111110",
1304 => "0000000000000001000000000100101100000000000000110101100000001",
1305 => "0000000000100011000000000000001100000001001010010101100000100",
1306 => "0000000001010001000000000000001100000000000001010101100000111",
1307 => "0000000000000001000000000000001100000000000000110101100001010",
1308 => "0000000000000001000000000000010100000000000000110101100001101",
1309 => "0000000000000001000000000000001100000000000001010101100010000",
1310 => "0000000000000001000000000000001100000000000000110101100010010",
1311 => "0000001010000010000000000000001100000000010010010101100010100",
1312 => "0000000000000001000000000000000100000000000000110101100010110",
1313 => "0000000000000001000000000000001100000000000000010101100011001",
1314 => "0000000000000001000000000010101100000000000000110101100011011",
1315 => "0000000000000001000000001010001000000000000000110101100011101",
1316 => "0000000000000001000000000000000100000000000000110101100100000",
1317 => "0000000000000001000000000000010100000000000000110101100100010",
1318 => "0000000000000001000000000000001100000000000010010101100100100",
1319 => "0000000000000001000000010000010000000000000000110101100100110",
1320 => "0000000000000001000000000000001100000000000000110101100101000",
1321 => "0000000000100001000000000000001100000000000001010101100101010",
1322 => "0000000000000001000000000000001100000000000000110101100101100",
1323 => "0000000100000010000000000000001100000000000000110101100101110",
1324 => "0000000000000011000000000000000100000000000000110101100110000",
1325 => "0000000000000001000000000000000100000000000000110101100110010",
1326 => "0000000000101011000000000000001100000000000000010101100110101",
1327 => "0000000000000001000000000000001100000000000000110101100111000",
1328 => "0000000000000001000000000000001100000000000000010101100111010",
1329 => "0000000000000001000000000000001100000000000000010101100111100",
1330 => "0000010000010101000000000000001100000000000000110101100111111",
1331 => "0000000000000001000000000001010100000000000001010101101000010",
1332 => "0000000000000001000000000000001100000000000000010101101000100",
1333 => "0000000000000001000000000000001100000000101010100101101000110",
1334 => "0000101010100100000000000000001100000000000000110101101001000",
1335 => "0000000000000001000000000000001100000000000000010101101001010",
1336 => "0000000000010001000000000000010100000000000000110101101001101",
1337 => "0000000000000001000000000000001100000000000001010101101010000",
1338 => "0000000000000001000000000000001100000000000000110101101010010",
1339 => "0000000000000101000000000000001100000000000000010101101010100",
1340 => "0000000000000001000000000000000100000000000000110101101010110",
1341 => "0000000000000001000000000010101100000000000000110101101011000",
1342 => "0000000000000001000000000000001100000000000000110101101011010",
1343 => "0000000000000001000000000000001100000000000000010101101011100",
1344 => "0000000000000001000000000000000100000000000000110101101011110",
1345 => "0000000000000101000000000000001100000000000000010101101100000",
1346 => "0000000000000001000000000000001100000000000000110101101100010",
1347 => "0000000000000001000000000000001100000001001001010101101100100",
1348 => "0000000000000001000000000000001100000000000000110101101100110",
1349 => "0000000000000011000000000000000100000010101010100101101101001",
1350 => "0000000000000001000000000000000100000000000000110101101101011",
1351 => "0000000000000001000000000000001100000000000000010101101101101",
1352 => "0000000000000001000000000000001100000000000000110101101101111",
1353 => "0000000000000011000000000000000100000000000000110101101110001",
1354 => "0000000000000001000000010010101000000000000000110101101110100",
1355 => "0000010100100000000000000000000100000000000000110101101110111",
1356 => "0000000000000011000000000001001100000000000000110101101111010",
1357 => "0000000000000001000000000000001100000000000000010101101111100",
1358 => "0000000000000101000000000000001100000000000000110101101111110",
1359 => "0000000000000001000000000000001100000000000000110101110000000",
1360 => "0000000000000001000000000000010100000000000000110101110000010",
1361 => "0000000000000001000000000000001100000000000000010101110000100",
1362 => "0000000000000001000000000000001100000000000101000101110000110",
1363 => "0000000000000001000000000001001100000000000000010101110001000",
1364 => "0000000000000001000000000000001100000000000000110101110001010",
1365 => "0000000000000001000000001000100100000000000000110101110001100",
1366 => "0000000000000001000000000000001100000000000000110101110001110",
1367 => "0000000000010011000000001000100000000000000000110101110010000",
1368 => "0000000001010001000000000000001100000000000000010101110010010",
1369 => "0000000000000001000000000000000100000000000000110101110010100",
1370 => "0000000000000001000000000000001100000000000000010101110010110",
1371 => "0000000000000001000000000000000100000000000000010101110011001",
1372 => "0000000000000001000000000000000100000000000000110101110011100",
1373 => "0000000000000001000000000000001100000000000100010101110011111",
1374 => "0000000000000001000000000000001100000000000000110101110100001",
1375 => "0000000000000001000000000000001100000000000100010101110100011",
1376 => "0000000000000001000000000000001100000000000000010101110100101",
1377 => "0000000000000001000000000000010100000000000010000101110100111",
1378 => "0000000000001011000000000000001100000010001010010101110101010",
1379 => "0000000000000001000000101000010000000000000000110101110101100",
1380 => "0000000000000001000000000000001100000000000000010101110101110",
1381 => "0000000000000001000000000000001100000000000000110101110110000",
1382 => "0000000000000001000000000000001100000000000100000101110110010",
1383 => "0000000000000001000000000000001100000000010010010101110110100",
1384 => "0000000000000001000000000000001100000000000000110101110110110",
1385 => "0000000000000001000000000000000100000000000000110101110111000",
1386 => "0000000000000001000000000000001100000000000000110101110111010",
1387 => "0000001000100010000000000000001100000000000000010101110111100",
1388 => "0000000000000001000000000000000100000000000000110101110111110",
1389 => "0000000000000001000000000000001100000001000101010101111000000",
1390 => "0000000000000001000000000000001100000000000000110101111000011",
1391 => "0000000000000001000000000000000100000000000000110101111000110",
1392 => "0000000000000001000000000000000100000000000000110101111001000",
1393 => "0000000000001001000000000000000100000000000000110101111001010",
1394 => "0000000000000001000000000000000100000000000000110101111001100",
1395 => "0000000000000001000000000000010100000000000000010101111001110",
1396 => "0000000000000001000000000000000100000000000000110101111010000",
1397 => "0000000000000001000000000000001100000000010010010101111010010",
1398 => "0000000000000001000000000000001100000000000000110101111010100",
1399 => "0000000000000001000000000000001100000000001000010101111010110",
1400 => "0000000000001011000000000001001100000000000000110101111011000",
1401 => "0000000000010101000000000000100100000000000000110101111011010",
1402 => "0000000000000001000000000000001100000000000000010101111011100",
1403 => "0000000100100001000000000000100100000000000000110101111011110",
1404 => "0000000000000001000000000000001100000000000000010101111100000",
1405 => "0000000000001001000000000000001100000000000000010101111100010",
1406 => "0000000000000001000000000000001100000000000000010101111100100",
1407 => "0000000000000001000000000001010100000000000000110101111100110",
1408 => "0000000000000001000000000000100100000000000000110101111101001",
1409 => "0000000000000001000000000000000100000000000000110101111101100",
1410 => "0000010000100101000000000000001100000000000010010101111101110",
1411 => "0000000000000001000000000000001100000000000000010101111110000",
1412 => "0000000000100100000000000000001100000000001000110101111110011",
1413 => "0000000000000000000000000000001100000000000000010101111110101",
1414 => "0000000000000001000000000000001100000000000000010101111110111",
1415 => "0000000010000100000000000000100100000000000000110101111111001",
1416 => "0000000000000001000000000000001100000000000000010101111111011",
1417 => "0000000000000001000000000000001100000000000000110101111111101",
1418 => "0000000000000011000000001000101000000000000000110101111111111",
1419 => "0000000000000001000000000000001100000000000000010110000000001",
1420 => "0000000000000001000000000000001100000000000000010110000000011",
1421 => "0000000000000001000000000000001100000000000000010110000000101",
1422 => "0000000000000001000000000000001100000000000010110110000000111",
1423 => "0000000000000001000000000010010000000000000000110110000001001",
1424 => "0000000000000001000000000000001100000000000000110110000001011",
1425 => "0000000000000001000000000000000100000000000000110110000001110",
1426 => "0000000000000001000000000000001100000000000000010110000010000",
1427 => "0000000000000001000000000000000100000000000000110110000010010",
1428 => "0000000000000001000000000000001100000000000100110110000010101",
1429 => "0000000000000001000000000000010100000000000000110110000010111",
1430 => "0000000000000001000000000000001100000000000000010110000011001",
1431 => "0000000000001001000000000001000100000000000000110110000011011",
1432 => "0000000000000001000000000000001100000000000001010110000011101",
1433 => "0000000000000001000000000000001100000000000000010110000011111",
1434 => "0000000000000001000000000000010100000000000000110110000100001",
1435 => "0000000000000001000000000000001100000000000000110110000100011",
1436 => "0000000000000101000000000100001100000000000000110110000100101",
1437 => "0000000000000001000000000000001100000000000000110110000100111",
1438 => "0000000000000001000000000000000100000000000000110110000101001",
1439 => "0000000000000001000000000000010100000000000000110110000101011",
1440 => "0000000000000001000000000001010000000000000000010110000101101",
1441 => "0000000000000001000000000000001100000000000000010110000101111",
1442 => "0000000000000001000000000000001100000000000001010110000110001",
1443 => "0000000000000001000000000000001100000000000000110110000110011",
1444 => "0000000010100001000000000000000000000001000010110110000110101",
1445 => "0000000000001001000000000000001100000000000000110110000110111",
1446 => "0000000000000001000000000001001100000000000000110110000111001",
1447 => "0000000000000001000000000000010100000000000000110110000111011",
1448 => "0000000000000001000000000000001100000000000010110110000111101",
1449 => "0000000000001011000000000000001100000000000000110110001000000",
1450 => "0000000000000011000000000001010100000000000000110110001000010",
1451 => "0000000000000001000000000000001100000000000000010110001000100",
1452 => "0000000000000001000000000000100100000000000000110110001000111",
1453 => "0000000000000001000000000000001100000000000010010110001001001",
1454 => "0000000000000001000000000000001100000000000000010110001001011",
1455 => "0000000000000001000000000000000100000000000000110110001001101",
1456 => "0000000000000001000000000010101100000000000000110110001001111",
1457 => "0000000000000001000001010010000100000000000000110110001010001",
1458 => "0000000000000001000000000000001100000000000000010110001010011",
1459 => "0000000000000001000000101000100000000000000000110110001010101",
1460 => "0000000000000001000000000000001100000000000000110110001011000",
1461 => "0000000000000001000000000000001100000000000000110110001011010",
1462 => "0000000000000001000000000000001100000000100000010110001011100",
1463 => "0000000000000001000000000000000100000000000000110110001011110",
1464 => "0000000100001001000000000000001100000000000000010110001100000",
1465 => "0000000000000001000000000000001000000000000000110110001100010",
1466 => "0000000001000000000000000000001100000001010010100110001100100",
1467 => "0000000000000001000000000000001100000000000000110110001100110",
1468 => "0000000000000001000000000000000100000000000000110110001101000",
1469 => "0000000000000101000000000000001100000000001001010110001101011",
1470 => "0000000000000001000000000000001100000000100000000110001101110",
1471 => "0000000000000001000000000000001100000000000000110110001110001",
1472 => "0000000000010001000000000000000100000000000000110110001110011",
1473 => "0000000000000001000000000000000100000000000000110110001110110",
1474 => "0000000000000001000000001000000000000000000000110110001111000",
1475 => "0000000000001001000000000000001100000000000000110110001111010",
1476 => "0000000000000001000000100001001000000000000100010110001111100",
1477 => "0000000000000011000000000000001100000000000000110110001111110",
1478 => "0000000100010100000000000000000100000000000000110110010000000",
1479 => "0000000000000001000000000000000100000000000000110110010000010",
1480 => "0000000000000101000000000000000100000000000000110110010000100",
1481 => "0000000000001011000000000000001100000000000000110110010000110",
1482 => "0000000001000001000000000000101100000000000000110110010001000",
1483 => "0000000000000001000000000000001100000000000000110110010001011",
1484 => "0000000000000001000000000000100100000000000000110110010001110",
1485 => "0000000000000101000000000000001100000000000000110110010010001",
1486 => "0000000000000001000000000000000100000000000000110110010010100",
1487 => "0000000000000001000000000000001100000000000010110110010010110",
1488 => "0000000000000001000000000000000100000000000000110110010011001",
1489 => "0000000000000001000000000000000100000000000000110110010011100",
1490 => "0000000000001001000000000000001100101000000000000110010011111",
1491 => "0000000000001011000000000000001100000001010101010110010100010",
1492 => "0000000000000001000000000000001100000000000000110110010100101",
1493 => "0000000000000001000000000000001100000000010101010110010100111",
1494 => "0000000000000011000000000000000100000000000000110110010101010",
1495 => "0000000000000001000000000000001100000000000000110110010101100",
1496 => "0000000000000001000000000000000100000000000000010110010101110",
1497 => "0000000000000001000000100101001000000000000000110110010110001",
1498 => "0000000000000001000000000000010100000100010101000110010110100",
1499 => "0000000000000101000000000000001100000000000000010110010110110",
1500 => "0000000000000001000000000000101100000000000010010110010111000",
1501 => "0000000000000101000000000000001100000000000000110110010111011",
1502 => "0000000000000011000000000000001100000000000000110110010111101",
1503 => "0000000000000001000000000000000100000000000000110110011000000",
1504 => "0000000000000001000000000000001100000000000000010110011000011",
1505 => "0000000000000001000000000000000100000000000000110110011000110",
1506 => "0000000000000001000000000000001100000000000000110110011001001",
1507 => "0000001000000100000000000000001100000000000000110110011001011",
1508 => "0000000000000001000000000000001100000000000000110110011001101",
1509 => "0000000000000001000000000000001100000000000000110110011001111",
1510 => "0000000000000001000000000000000100000000000000010110011010001",
1511 => "0000000000101001000000000000001100000000000000110110011010100",
1512 => "0000000000000001000000000000001100000000000000010110011010111",
1513 => "0000000000000001000000000000001100000000000000110110011011001",
1514 => "0000000000000001000000000000001100000000000000010110011011100",
1515 => "0000000000000001000000000000000100000000000000110110011011110",
1516 => "0000000000000001000000000000001100000000010000110110011100001",
1517 => "0000000000000001000000000000001100000000000000010110011100011",
1518 => "0000000000000101000000000000001100000000000000110110011100101",
1519 => "0000000000000001000000000000000100000000000000110110011100111",
1520 => "0000000000000001000000000000001100000000000000010110011101001",
1521 => "0000000000000001000000000000001100000000000000010110011101100",
1522 => "0000000000000001000000000000001100000000000100010110011101111",
1523 => "0000000000000011000000000000001100000000000000010110011110001",
1524 => "0000000000001001000000000101001100000000000000110110011110011",
1525 => "0000000000000001000000000000000100000000000000110110011110101",
1526 => "0000000000000001000000000000010100000000000000110110011110111",
1527 => "0000000000000001000000000000001100000000000000110110011111001",
1528 => "0000000000000011000000001000000000000000000000110110011111011",
1529 => "0000000000000011000000000000001100000000000000110110011111101",
1530 => "0000000000000001000000000000101100000000000000010110011111111",
1531 => "0000000000000101000000000000001100000000000000110110100000010",
1532 => "0000000000000001000000000010100100000000000000010110100000100",
1533 => "0000000000001011000000000000000100000000000000110110100000110",
1534 => "0000000000000001000001000010001000000000010001010110100001000",
1535 => "0000000000000001000000000000001100000000000000110110100001010",
1536 => "0000000000000001000000000000001100000000000001010110100001100",
1537 => "0000000000100011000000000000001100000000000000110110100001110",
1538 => "0000000000000011000000000000000100000000000000010110100010000",
1539 => "0000000000000011000000000000001100000000000000110110100010010",
1540 => "0000000010101001000000000100101100000000000000110110100010100",
1541 => "0000000000001011000000000000001100000000000000110110100010110",
1542 => "0000000000000001000000000000001100000000000000010110100011000",
1543 => "0000000000000001000000000000001100000000000000110110100011011",
1544 => "0000000000000001000000000000000100000000000000010110100011101",
1545 => "0000000000000001000000000000001100000000000000110110100011111",
1546 => "0000000000000001000000000000001100000000000000010110100100001",
1547 => "0000000000000001000000000000001100000000000000110110100100011",
1548 => "0000000000000001000000000000101100000000000000110110100100101",
1549 => "0000000000000001000000000000001100000001000010000110100101000",
1550 => "0000000000000001000000000000001100000000000000110110100101010",
1551 => "0000000000000001000000000000000100000000000000110110100101100",
1552 => "0000000000001011000000000000000100000000000001010110100101110",
1553 => "0000000000000001000000000000000100000000000000110110100110000",
1554 => "0000000000000001000000000000001100000000000000010110100110010",
1555 => "0000000000000001000000000000001100000000010001010110100110100",
1556 => "0000000000001001000000000000001100000000010000110110100110110",
1557 => "0000010000010011000000000010001100000000000000110110100111001",
1558 => "0000000000000001000000000000101100000000010100000110100111011",
1559 => "0000000000000001000000000000001100000000100000010110100111101",
1560 => "0000000000000001000000000000001100000000000000110110100111111",
1561 => "0000000000000001000000000000001100000000000001010110101000001",
1562 => "0000000100000100000000000000001100000000000000010110101000011",
1563 => "0000000000000001000000000000001100000000000001010110101000101",
1564 => "0000000000000001000000000000001100000010000001000110101000111",
1565 => "0000000101001000000000000000001100000000000000010110101001001",
1566 => "0000000000000001000000000000001100000000000000010110101001100",
1567 => "0000000000000001000000000000001100000000000000010110101001111",
1568 => "0000000000001011000000000000001100000000000000110110101010001",
1569 => "0000000000000001000000000010101100000000001010000110101010011",
1570 => "0000000000000001000000000000001100000000000000110110101010101",
1571 => "0000000000000001000000000000001100000000000000010110101010111",
1572 => "0000000000000001000000100000001100000000000000110110101011010",
1573 => "0000000000000001000000000000001100000000000000010110101011100",
1574 => "0000000000000001000000000000001100000000000101010110101011110",
1575 => "0000000000000001000000001000101100000000000000110110101100000",
1576 => "0000000000100101000000000000001100000000000000010110101100010",
1577 => "0000000000000001000000000000001100000000000001010110101100101",
1578 => "0000000000000001000000000000001100000000000000110110101101000",
1579 => "0000000000000001000000001010101000000000000000110110101101010",
1580 => "0000000000000001000000010100000100000000000000110110101101100",
1581 => "0000000000000001000000000000001100000001000100000110101101110",
1582 => "0000000000000001000000000000001100000000000000010110101110000",
1583 => "0000000000000001000000000000001100000000000000010110101110010",
1584 => "0000000000000001000000000000000100000000000000110110101110101",
1585 => "0000000000000001000000000000001100000000000010010110101110111",
1586 => "0000000100000000000000000000001100000000000000110110101111001",
1587 => "0000000100100010000000000000001100000000001000010110101111011",
1588 => "0000000000000001000000000000001100000000000000110110101111101",
1589 => "0000000000000001000000000000001100000000100101000110101111111",
1590 => "0000000000000001000000000000001100000000000000010110110000001",
1591 => "0000000000000001000000000000001100000000010000010110110000011",
1592 => "0000000000000001000000000000001100000000000000010110110000101",
1593 => "0000000000000001000000000000001100000000000100010110110000111",
1594 => "0000000000000001000000000000000100000000000000110110110001001",
1595 => "0000000000000011000000000000001100000000000000110110110001011",
1596 => "0000000000000001000000000000001100000000000010010110110001101",
1597 => "0000000000000001000000000000001100000000000000110110110010000",
1598 => "0000000000000001000000000000001100000000000000110110110010010",
1599 => "0000000000000001000000000000001100000000000000010110110010100",
1600 => "0000000000001001000000000000001100000000100100100110110010110",
1601 => "0000000000101001000000000000001100000000000000110110110011000",
1602 => "0000000000000011000000000000001100000000000000110110110011010",
1603 => "0000000000000001000000000000000100000000000000010110110011100",
1604 => "0000001010000101000000000000001100000000000000110110110011110",
1605 => "0000000000000011000000000000001100000000000000010110110100000",
1606 => "0000000000000001000000000000001100000000000000010110110100011",
1607 => "0000000000000001000000000000001100000000000000010110110100101",
1608 => "0000000000000001000000000000000100000000000000110110110101000",
1609 => "0000000000000101000000000000001100000000010000010110110101010",
1610 => "0000000000000001000000000000000100000000000000110110110101100",
1611 => "0000000000000001000000010100101000000000000000110110110101111",
1612 => "0000000000000001000000000000001100000000000000110110110110001",
1613 => "0000000000000001000000000000001100000000000001010110110110100",
1614 => "0000000000010101000000000000001100000000000000010110110110110",
1615 => "0000000000000001000000000000101100000000000000110110110111000",
1616 => "0000000000000001000000000000001100000000000101000110110111010",
1617 => "0000000000000001000000000000000100000000001010010110110111100",
1618 => "0000000000000001000000000100001100000000000000110110110111110",
1619 => "0000000000000001000000001010000100000000000100010110111000000",
1620 => "0000000000000001000000000000001100000000000010010110111000010",
1621 => "0000000000000001000000000000001100000000101010010110111000100",
1622 => "0000100100001010000000000000001100000000000000110110111000110",
1623 => "0000000000100011000000000000001100000000000000010110111001000",
1624 => "0000000000000011000000000000001100000000000000110110111001010",
1625 => "0000000000010000000000000000001100000000000000010110111001100",
1626 => "0000000000001001000000000000001100000010001010010110111001110",
1627 => "0000000000000001000000000000000100000000000000110110111010000",
1628 => "0000000000000001000000000000001100000001010010100110111010010",
1629 => "0000000000000001000000000000001100000000000000110110111010100",
1630 => "0000000000000001000000000000001100000000000000110110111010110",
1631 => "0000000000000001000000000000001100000000000000010110111011000",
1632 => "0000000000000001000000000000001100000000000000110110111011010",
1633 => "0000000000000001000000101000010000000000000001010110111011100",
1634 => "0000000000000001000000010101001100000000000000110110111011110",
1635 => "0000000000000001000000000000001100000000000010110110111100000",
1636 => "0000000000001001000000000000001100000000000000010110111100010",
1637 => "0000000000000001000000001001000000000000000000110110111100100",
1638 => "0000000000000001000000000000001100000000000000110110111100110",
1639 => "0000000000000001000000000000001100000000010100010110111101000",
1640 => "0000000000000001000000000000000100000000000000110110111101010",
1641 => "0000000000000001000000000000000100000000000000110110111101100",
1642 => "0000000000000001000000000000001100000000000000110110111101110",
1643 => "0000000000000001000000000000001100000000100100100110111110000",
1644 => "0000000000000001000000000000001100000000000001000110111110010",
1645 => "0000000000000001000000000000001100000000000001010110111110100",
1646 => "0000000010001001000000000000000100000000000000110110111110110",
1647 => "0000000000000001000000000000001100000000000010010110111111000",
1648 => "0000000000000001000000000000001100000000000010110110111111010",
1649 => "0000000000000001000000000000000100000000000000110110111111101",
1650 => "0000000000000011000000000000001100000001010101010110111111111",
1651 => "0000000000000001000000000000001100000000000010010111000000001",
1652 => "0000000000100101000000000001001000000000000000110111000000100",
1653 => "0000000000000101000000000000001100000010001010100111000000111",
1654 => "0000000000101001000000000000001100000000000000010111000001010",
1655 => "0000000000000001000000000000000100000000000000110111000001100",
1656 => "0000000010000101000000000000001100000000000000110111000001110",
1657 => "0000000000000011000000000000001100000000000000010111000010000",
1658 => "0000010100000100000000000000001100000000000000110111000010011",
1659 => "0000000000000001000000000000000100000000000000110111000010110",
1660 => "0000000000000001000000000000001100000000000001010111000011000",
1661 => "0000000000000001000000000000001100000000010010110111000011011",
1662 => "0000000000000001000000000000001100000000000000110111000011101",
1663 => "0000000000000101000000000000001100000000000000010111000011111",
1664 => "0000000000000001000000000000001100000000000000010111000100001",
1665 => "0000000000000001000000000000000100000000000000110111000100011",
1666 => "0000000000000001000000000000001100000000000001010111000100101",
1667 => "0000000000000001000000000000001100000001000000000111000100111",
1668 => "0000000000000001000000000000001100000000000010110111000101001",
1669 => "0000000000000001000000000000000100000000000000110111000101100",
1670 => "0000000000000001000000000100101100000000000000110111000101111",
1671 => "0000000000000001000000000000000100000000000010100111000110001",
1672 => "0000000000000011000000000000001100000000000000010111000110011",
1673 => "0000000000000001000000000000001100000000000000110111000110101",
1674 => "0000000000000001000000000000001100000000000010010111000110111",
1675 => "0000000000000011000000000001001000000000001010010111000111001",
1676 => "0000000000000001000000000001000100000000000000110111000111011",
1677 => "0000000000000001000000000000010100000000000000110111000111101",
1678 => "0000000000000001000000000000001100000000000000010111001000000",
1679 => "0000000000000001000000000000000100000000000000110111001000010",
1680 => "0000000000000001000000000000001100000000000000110111001000100",
1681 => "0000000000001001000000000000001100000010010010010111001000111",
1682 => "0000000000000001000000000000010100000000000000110111001001001",
1683 => "0000000000000001000000000001010100000000000000110111001001011",
1684 => "0000001010000101000000000000001100000000010000110111001001110",
1685 => "0000000000000001000000000000001100000000100100100111001010001",
1686 => "0000000000000001000000000000001100000000100010110111001010100",
1687 => "0000000000000001000000001001000100000000000000110111001010110",
1688 => "0000000000000001000000000000000100000000000000110111001011000",
1689 => "0000000000000001000000000000001100000000000100010111001011010",
1690 => "0000000000000001000000000000001100000000000000110111001011100",
1691 => "0000000000000001000000000010001000000000001001010111001011110",
1692 => "0000000000000001000000000000001100000000000000110111001100000",
1693 => "0000000000100001000000000001010000000000000000110111001100010",
1694 => "0000000000000001000000000000000100000000000000110111001100100",
1695 => "0000000101000010000000000000001100000000000000110111001100110",
1696 => "0000000000000011000000000000001100000000000000110111001101000",
1697 => "0000000000001001000000000000000100000000000000110111001101010",
1698 => "0000000100010100000000000000001100000000000001010111001101100",
1699 => "0000000000000001000000000000000100000000001000010111001101110",
1700 => "0000000000000001000000000010100100000000000000110111001110000",
1701 => "0000000000000001000000000000001100000000000000110111001110010",
1702 => "0000000000000001000000000000000100000000000000110111001110100",
1703 => "0000000000000001000000001000101100000000000000010111001110111",
1704 => "0000000000000001000000000000010100000000000000110111001111001",
1705 => "0000000010000101000000001010001000000000000000110111001111011",
1706 => "0000000000000001000000000000001100000000000000110111001111101",
1707 => "0000000010100001000000000000001100000000000001010111001111111",
1708 => "0000000000000001000000000000001100000000000000110111010000001",
1709 => "0000000000000011000000000000001100000000000101010111010000011",
1710 => "0000000010000101000000000000001100000000000000010111010000101",
1711 => "0000000000000011000000000000000100000000000011110111010000111",
1712 => "0000000000000001000000000000001100000000000000110111010001001",
1713 => "0000000000000001000000000101001100000000000000110111010001011",
1714 => "0000000000000101000000000000001100000000000000110111010001110",
1715 => "0000000000000011000000000000000100000000000000110111010010000",
1716 => "0000000000000001000000000000001100000000000000110111010010010",
1717 => "0000000010000101000000000000100100000000000000110111010010100",
1718 => "0000000000000001000000000000101100000000000000110111010010110",
1719 => "0000000000000001000000000000001100000000001000010111010011000",
1720 => "0000000000000001000000000100000100000000000000110111010011010",
1721 => "0000000000000001000000000000001100000000000010010111010011101",
1722 => "0000000001000100000000000000001100000000000000010111010011111",
1723 => "0000000000000001000000000000101100000000000000110111010100001",
1724 => "0000000000000001000000000000001100000000000000110111010100011",
1725 => "0000000000000001000000000000000100000000000000110111010100101",
1726 => "0000000000000001000000000000001100000000000000110111010100111",
1727 => "0000000000000001000000000010001000000000000000010111010101010",
1728 => "0000000000000001000000000001000100000000000000110111010101100",
1729 => "0000000001001001000000000000001100000000000001010111010101110",
1730 => "0000000000000001000000000000001100000000000000010111010110000",
1731 => "0000000001010011000000000000001100000000000010010111010110010",
1732 => "0000100000010101000000000000001100000000000000010111010110100",
1733 => "0000000101010010000000000000000100000000000000110111010110110",
1734 => "0000001000000001000000000000001100000000000000110111010111000",
1735 => "0000000000000001000000000000000100000000000000110111010111010",
1736 => "0000000000000001000000000000001100000000010000010111010111100",
1737 => "0000000000000001000000000000000100000000000000110111010111110",
1738 => "0000000000100011000000000000001100000000001000010111011000000",
1739 => "0000000000000001000000000000001100000000000000110111011000010",
1740 => "0000000000000001000000000000001100000000000000010111011000100",
1741 => "0000000000000001000000000000000100000000000000110111011000110",
1742 => "0000000000000001000000000000001100000000000000010111011001000",
1743 => "0000000000000001000000000000001100000000000000110111011001010",
1744 => "0000000000000101000000000000001100000000000010010111011001100",
1745 => "0000000000000001000000000000001100000001000100100111011001110",
1746 => "0000000000000101000000000000000100000000000000110111011010000",
1747 => "0000000000000001000000000000000100000000000000110111011010010",
1748 => "0000000000101011000000000000001100000000000000010111011010100",
1749 => "0000000000000011000000000000001100000000000000010111011010110",
1750 => "0000000000000001000000000000001100000000100100100111011011000",
1751 => "0000000000100101000000000000001100000000000000110111011011010",
1752 => "0000000000000001000000000001000100000000000000110111011011101",
1753 => "0000000000000001000000000000001100000000000000000111011011111",
1754 => "0000000000000001000000000000001100000000101010000111011100001",
1755 => "0000000000000001000000000000001100000000000000010111011100011",
1756 => "0000000000000001000000000000000100000000000000110111011100101",
1757 => "0000000000000011000000000000001100000000000000110111011100111",
1758 => "0000000000000001000000000000001100000000000001010111011101001",
1759 => "0000000000000011000000000000001100000000010000010111011101011",
1760 => "0000000000001001000000000000001100000001001010000111011101101",
1761 => "0000000000000001000000000000001100000000000000110111011101111",
1762 => "0000000000000001000000000000010100000000000000110111011110001",
1763 => "0000000000000001000000000000001100000000000000110111011110011",
1764 => "0000000000000011000000000001000100000000000000010111011110110",
1765 => "0000000000000001000000000000000100000000000000110111011111001",
1766 => "0000000000100101000000000000001100000000000010010111011111011",
1767 => "0000000000000001000000000000001100000000000000110111011111110",
1768 => "0000000000000001000000000001010100000000000000110111100000000",
1769 => "0000000000000101000000000000000100000000000000110111100000011",
1770 => "0000000000000011000000000000001100000001010100000111100000110",
1771 => "0000000000000001000000000000101100000000000000110111100001000",
1772 => "0000000001010011000000000000001100000001001010010111100001010",
1773 => "0000000000000001000000000000001100000000000000110111100001100",
1774 => "0000000000000001000000000000001100000000000000010111100001110",
1775 => "0000000000001011000000000000101100000000000000110111100010000",
1776 => "0000000000000001000000000000001100000000000001010111100010010",
1777 => "0000000000000101000000000010010100000000000000110111100010100",
1778 => "0000000000000001000000000000001100000000000000010111100010110",
1779 => "0000000000001001000000000000001100000000100001010111100011000",
1780 => "0000000000000001000000000000001100000000100100000111100011010",
1781 => "0000000000000101000000000000001100000000000100110111100011100",
1782 => "0000000000100011000000000000001100000000000000010111100011110",
1783 => "0000000000000001000000000000001100000000000000110111100100000",
1784 => "0000000000000001000000001010101000000000000000110111100100010",
1785 => "0000000000000001000000000000001100000000000000110111100100100",
1786 => "0000000000000011000000000000000100000000000000110111100100110",
1787 => "0000000000000001000000000000100100000000000000110111100101001",
1788 => "0000000000000001000000000000100100000000000000110111100101011",
1789 => "0000000000000001000000000000001100000000000000110111100101101",
1790 => "0000000000000001000000001001000100000000000000110111100110000",
1791 => "0000000000000001000000000000000100000000000000110111100110010",
1792 => "0000000000000001000000000000001100000000000000010111100110101",
1793 => "0000000000001011000000000000001100000000000000010111100110111",
1794 => "0000000000000001000000000000001100000000000000010111100111001",
1795 => "0000000001000011000000000000001100000000000000110111100111011",
1796 => "0000000000000001000000000000001100000001000001000111100111101",
1797 => "0000000000000011000000000000001100000000000000010111100111111",
1798 => "0000000000000001000000000000000100000000000000110111101000001",
1799 => "0000000000000001000000000000001100000000001000100111101000011",
1800 => "0000000000000001000000000001010100000000000000010111101000101",
1801 => "0000000000000001000000000000001100000000000000110111101001000",
1802 => "0000000000000001000000000000001100000000000001010111101001010",
1803 => "0000000000000001000000000000001100000000000000010111101001100",
1804 => "0000000000000001000000000000001100000000000000110111101001110",
1805 => "0000000000000001000000000000001100000000001010010111101010000",
1806 => "0000000000000001000000000000001100000000000000010111101010011",
1807 => "0000000000010001000000000000001100000000010000000111101010101",
1808 => "0000000000000001000000000000001100000000000000010111101010111",
1809 => "0000000000000001000000000000001100000000000000110111101011001",
1810 => "0000000000010011000000000000000100000000000000010111101011011",
1811 => "0000000000000011000000000000001100000000000000010111101011110",
1812 => "0000000000000001000000000000000100000000000000110111101100000",
1813 => "0000000000011011000000000000001100000000000000110111101100010",
1814 => "0000000000000001000000000000001100000000101000100111101100101",
1815 => "0000000000000101000000000000001100000000000000010111101100111",
1816 => "0000000000000001000000000000000100000000000000110111101101001",
1817 => "0000000000000011000000000000000100000000000000110111101101100",
1818 => "0000000001000011000000000000101100000000000000110111101101110",
1819 => "0000000000000001000000000000001100000000000000110111101110000",
1820 => "0000000000000001000000000000010100000000010101010111101110010",
1821 => "0000000000000101000000000000001100000000000010010111101110101",
1822 => "0000000000000001000000010100000100000000000000110111101111000",
1823 => "0000000000000001000000000000001100000000000000110111101111010",
1824 => "0000000000000011000000000000001100000010000001000111101111100",
1825 => "0000000000000001000000000000001100000000000001010111101111110",
1826 => "0000000001000011000000001001000000000000000000110111110000000",
1827 => "0000000000000101000000000000001100000000000000010111110000010",
1828 => "0000000000010101000000000000001100000000000000010111110000100",
1829 => "0000000100000101000000000000000100000000000000110111110000110",
1830 => "0000000000010001000000000000001100000000000000110111110001000",
1831 => "0000000000000001000000000000001100000000000000110111110001011",
1832 => "0000000000000001000000000000001100000000101000100111110001101",
1833 => "0000000000000001000000000000000100000000000000110111110001111",
1834 => "0000000000000001000000000000001100000000000001010111110010010",
1835 => "0000000000000001000000000000001100000000000000010111110010100",
1836 => "0000000000000001000000000000001100000000100101010111110010110",
1837 => "0000000000000001000000000000001100000001000100100111110011000",
1838 => "0000000000101011000000000000100100000000000000010111110011011",
1839 => "0000000000000001000000000000001100000000000000110111110011110",
1840 => "0000000010010101000000000001000100000000000000110111110100000",
1841 => "0000000010101001000000000000001100000000000000110111110100011",
1842 => "0000000100000001000000000000001100000000000000110111110100110",
1843 => "0000000000000001000000000000001100000000000000110111110101000",
1844 => "0000000000000001000000000000001100000000000000010111110101010",
1845 => "0000000000000001000000000000000100000000000000110111110101100",
1846 => "0000000000000001000000000000001100000000000000010111110101110",
1847 => "0000000000000001000000000000001100000000000000110111110110000",
1848 => "0000000000000001000000000001010100000000000000110111110110010",
1849 => "0000000000000001000000000000000100000000000000110111110110100",
1850 => "0000000000000001000000000000001100000000000010010111110110110",
1851 => "0000000000000001000000000000001100000000000001010111110111000",
1852 => "0000000000000001000000000100101100000000000000110111110111010",
1853 => "0000000000000001000000000000001100000000000000110111110111100",
1854 => "0000000001000101000000000000001100000001000000010111110111110",
1855 => "0000000100000101000000000000001100000000000100010111111000000",
1856 => "0000000000000001000000000000001100000000101000110111111000010",
1857 => "0000000000000001000000000000000100000000000000110111111000100",
1858 => "0000000000010001000000000000010100000000000000110111111000110",
1859 => "0000000000000001000000000000001100000000000000110111111001000",
1860 => "0000000000000001000000000000000100000000000000110111111001010",
1861 => "0000000000001001000000000000001100000000001010010111111001100",
1862 => "0000000000000001000000000000001100000000000010110111111001110",
1863 => "0000000000000001000000000000010100000000000000110111111010001",
1864 => "0000000000000001000000000000001100000000000000010111111010011",
1865 => "0000000000000001000000000000001100000000000000110111111010101",
1866 => "0000000000000001000000000000001100000000101010100111111010111",
1867 => "0000000000000001000000000000001100000100100000100111111011001",
1868 => "0000000000000001000000000000100100000000001001000111111011011",
1869 => "0000000000000001000000000000001100000000000000110111111011101",
1870 => "0000101010001000000000000000001100000010001010000111111011111",
1871 => "0000000000000001000000000000001100000000000000110111111100001",
1872 => "0000000000000001000000000000001100000000000000010111111100011",
1873 => "0000000000000001000000000000001100000000100000000111111100101",
1874 => "0000000000000001000000000000001100000000000000010111111100111",
1875 => "0000000000000001000000000000010100000000000000110111111101010",
1876 => "0000000000000001000000000000001100000000000000010111111101100",
1877 => "0000000000000001000000000000001100000000000000110111111101110",
1878 => "0000000000000011000000000000001100000000000000010111111110000",
1879 => "0000000000000001000000000001010100000000000000110111111110010",
1880 => "0000000000000001000000000000001100000000000001010111111110100",
1881 => "0000000000000001000000000000001100000000000000110111111110111",
1882 => "0000000001010101000000000100001100000000000000110111111111001",
1883 => "0000000000000001000000000000001100000000000000110111111111011",
1884 => "0000000000000011000000001010101000000000000000110111111111110",
1885 => "0000100000100011000000000000001100000000000000111000000000001",
1886 => "0000000000000101000000000000000100000000000000011000000000011",
1887 => "0000000000000001000000000000001100000000000000111000000000101",
1888 => "0000000000000001000000010010010100000000000000111000000000111",
1889 => "0000000000000001000000000000000100000000000000111000000001001",
1890 => "0000000000000101000000000000010100000000000000011000000001011",
1891 => "0000000000000001000000000000001100000000000000111000000001101",
1892 => "0000000000000001000000001010001100000000000001011000000001111",
1893 => "0000000000000001000000000000000100000000000000111000000010010",
1894 => "0000000000000001000000000000001100000000000000111000000010101",
1895 => "0000000000000001000000000000001100000001010100101000000010111",
1896 => "0000000000000001000000000000001100000000000000111000000011001",
1897 => "0000000000000001000000000000001100000000000000111000000011011",
1898 => "0000000000000001000000000000000100000000000010011000000011101",
1899 => "0000000000000001000000000000001100000000000000111000000011111",
1900 => "0000000001001001000000000000010100000000000000111000000100001",
1901 => "0000000000000001000000000000001100000000000000111000000100100",
1902 => "0000000000000001000000000100100100000000000000011000000100111",
1903 => "0000000001010001000000000010100100000000000000111000000101001",
1904 => "0000000000000001000000000000001100000000000000011000000101011",
1905 => "0000000000000001000000100000001000000000000000111000000101101",
1906 => "0000000000000001000000000000000100000000000000111000000101111",
1907 => "0000000000000001000000000000001100000000000000111000000110001",
1908 => "0000000000000001000000000000000100000000001000011000000110011",
1909 => "0000000000000101000000000000001100000000000000111000000110101",
1910 => "0000010000101000000000000001010100000000000000011000000110111",
1911 => "0000000000000101000000000000001100000000100000111000000111001",
1912 => "0000000010100101000000000000001100000000000000111000000111011",
1913 => "0000010101001000000000000000001100000000000000111000000111101",
1914 => "0000000000000001000000000000001100000000000000111000001000000",
1915 => "0000000000000001000000001010100100000000000000111000001000011",
1916 => "0000000000000001000000000000000100000000000000011000001000110",
1917 => "0000000000010101000000000000001100000000000010111000001001000",
1918 => "0000000000000001000000000000001100000000000000011000001001011",
1919 => "0000000000000001000000010000100000000000000000111000001001101",
1920 => "0000000000000011000000000000000100000000000000111000001001111",
1921 => "0000000000000001000000000000001100000000000000111000001010001",
1922 => "0000000000000001000000010100001000000000000000111000001010011",
1923 => "0000000000000001000000001000000100000000000000111000001010101",
1924 => "0000000000001001000000010001000000000000000000111000001010111",
1925 => "0000000000000001000000000000001100000000000001011000001011001",
1926 => "0000000000000001000000000000001100000000000000111000001011011",
1927 => "0000000000000011000000000000001100000000000100111000001011101",
1928 => "0000000000000011000000000000001100000000100100011000001011111",
1929 => "0000000000000001000000000000001100000000000000111000001100001",
1930 => "0000000000000001000000000000001100000000000000011000001100011",
1931 => "0000101010100000000000000000000100000000000000111000001100101",
1932 => "0000000000000001000000000000001100000000000000011000001100111",
1933 => "0000000000000101000000000000001100000000000000011000001101001",
1934 => "0000000000000011000000000000001100000000010100011000001101011",
1935 => "0000000000000001000000000000000100000000000000111000001101101",
1936 => "0000000000000001000000000101001100000000000000111000001101111",
1937 => "0000000000000001000000000000001100000000000010111000001110001",
1938 => "0000000000000001000000000001010100000000000000111000001110011",
1939 => "0000000000000001000000000000000100000000000000111000001110101",
1940 => "0000000000000001000000000000001100000000000000111000001110111",
1941 => "0000000000100011000000000000001100000000000000011000001111010",
1942 => "0000000000000001000000000000001100000000100001001000001111100",
1943 => "0000000000000001000000000000001100000000000000011000001111110",
1944 => "0000000000000001000000000100001100000000000000111000010000000",
1945 => "0000000000000001000000000000001100000000000000111000010000010",
1946 => "0000000000000001000000010100010100000000000000111000010000100",
1947 => "0000000000010001000000000000000100000000000000111000010000111",
1948 => "0000000000000001000000000000001100000000101010101000010001010",
1949 => "0000100100100100000000000000001100000000000000111000010001100",
1950 => "0000000000000001000000000000001100000000100000011000010001111",
1951 => "0000000000000001000000000000001100000000010001001000010010010",
1952 => "0000000000000001000000000000001100000000101001001000010010101",
1953 => "0000000000000001000000000000001100000000000000111000010010111",
1954 => "0000000000000001000000000100000100000000000000111000010011001",
1955 => "0000000000010011000000000000001100000000000000111000010011011",
1956 => "0000000000000001000000000000001100000000000000111000010011101",
1957 => "0000000000000001000000000000001100000000000000111000010100000",
1958 => "0000000000000001000000001010100100000000000000111000010100010",
1959 => "0000000000000001000000000000001100000000000000011000010100101",
1960 => "0000000000000011000000000000001100000000000000111000010100111",
1961 => "0000000000000001000000000000001100000000000000011000010101001",
1962 => "0000000000000001000000000000001100000000000001011000010101011",
1963 => "0000000000000001000000000000000100000000000000111000010101101",
1964 => "0000000000000001000000000000001100000000010010011000010110000",
1965 => "0000000000000001000000000100010100000000000000111000010110010",
1966 => "0000000000000001000000000000001100000000000000011000010110100",
1967 => "0000000000000001000000000000001100000000000000111000010110110",
1968 => "0000000000101001000000000000010100000000000001011000010111001",
1969 => "0000000001010011000000000000001100000000000001011000010111011",
1970 => "0000000000000001000000000000001100000000010100011000010111101",
1971 => "0000000000000011000000000000101100000000000000111000010111111",
1972 => "0000000000000001000000000000001100000000000000011000011000001",
1973 => "0000000000000001000000000000000100000000000000111000011000011",
1974 => "0000000000000001000000000001000100000000001010001000011000101",
1975 => "0000000000000001000000000000001100000000100100011000011000111",
1976 => "0000000000000001000000000000000100000000000010111000011001001",
1977 => "0000000000000001000000000000001100000000000000111000011001011",
1978 => "0000000000000001000000000010001100000000000000011000011001101",
1979 => "0000000000000001000000000000100100000000000000111000011010000",
1980 => "0000000000010011000000000010001100000000000000111000011010010",
1981 => "0000000000000001000000000000001100000000000000111000011010100",
1982 => "0000000000000001000000000000001100000000000000111000011010110",
1983 => "0000000000000001000000000000001100000000000000111000011011000",
1984 => "0000000000000001000000000000001100000000000000011000011011010",
1985 => "0000000000000001000000000000000100000000000000111000011011100",
1986 => "0000000000000001000000000000001100000000000000111000011011111",
1987 => "0000000000000001000000000000001100000000000000111000011100001",
1988 => "0000000000000001000000000000000100000000000101001000011100011",
1989 => "0000000000000001000000000000001100000000000000011000011100101",
1990 => "0000000000010011000000000000001100000000000000111000011100111",
1991 => "0000000000000001000000000000000100000000000000111000011101001",
1992 => "0000010000010000000000000001000000000000000100111000011101011",
1993 => "0000000000000001000000000000000100000000000000111000011101110",
1994 => "0000001010000000000000000000001100000000000000111000011110000",
1995 => "0000000000000001000000000000001100000000000000111000011110010",
1996 => "0000000000000001000000000000001100000000000001011000011110100",
1997 => "0000000000000001000000000000001100000000000000011000011110110",
1998 => "0000000000000001000000000000001100000000000010011000011111000",
1999 => "0000000000000001000000000000000100000000000000111000011111010",
2000 => "0000000100001011000000000000000100000000000000111000011111100",
2001 => "0000000000000001000000000000001100000000000000111000011111110",
2002 => "0000000000000001000000000000001100000000000000111000100000000",
2003 => "0000000000000001000000000000000100000000000000111000100000010",
2004 => "0000000000000001000000000010101100000000000000111000100000101",
2005 => "0000000000000001000000000000001100000000000000111000100001000",
2006 => "0000000000100000000000000000001100000000000000111000100001011",
2007 => "0000000000000001000000000000000100000000000000111000100001101",
2008 => "0000000000000001000000000000000100000000000000111000100001111",
2009 => "0000000000000001000000000000001100000000000000111000100010001",
2010 => "0000000000000001000000000000000100000000000000111000100010100",
2011 => "0000000000000001000000000000001100000000000000111000100010110",
2012 => "0000000101010000000000000000001100000000000000011000100011000",
2013 => "0000000000000001000000000001010100000000000000111000100011010",
2014 => "0000000000100101000000000010010100000000000000011000100011100",
2015 => "0000000000000001000000000000001100000000000000111000100011110",
2016 => "0000000000000001000000010101010100000000000000011000100100001",
2017 => "0000000000000001000000000000000100000000000000111000100100011",
2018 => "0000000000100101000000000000001100000000000000011000100100110",
2019 => "0000000000000001000000010001000100000000000000111000100101000",
2020 => "0000000000000001000000000000001100000000000100011000100101011",
2021 => "0000000000000001000000000000001100000000000010011000100101110",
2022 => "0000000000000001000000000000001100000000001001011000100110001",
2023 => "0000000000000001000000000000000100000000000000111000100110011",
2024 => "0000100010001010000000000010001100000000000000111000100110101",
2025 => "0000000000000001000000000000001100000000000000011000100110111",
2026 => "0000000000000001000000000000000100000000000000111000100111010",
2027 => "0000000000000001000000000000001100000000000000111000100111100",
2028 => "0000000000000001000000010010100000000000000000111000100111110",
2029 => "0000000000000001000000000001010100000000000000111000101000000",
2030 => "0000000000000001000000000000001100000000000100111000101000010",
2031 => "0000000000000001000000000000001100000000000010111000101000100",
2032 => "0000010000010010000000000010100100000000000000111000101000110",
2033 => "0000000000100011000000000000001100000000000010111000101001000",
2034 => "0000000000000001000000000000000100000000000000011000101001010",
2035 => "0000000000000001000000000000001100000000000010111000101001100",
2036 => "0000000000000001000000000000001100000000000000011000101001110",
2037 => "0000000000000001000000000000001100000000000000011000101010001",
2038 => "0000000100000011000000000000001100000001000010011000101010011",
2039 => "0000000000000001000000000000001100000000000000111000101010101",
2040 => "0000000000000001000000010000001000000000000000111000101011000",
2041 => "0000000000000001000000000000001100000000000000111000101011011",
2042 => "0000000000000101000000000000000100000000000000011000101011110",
2043 => "0000000000000001000000000000000100000000000000111000101100001",
2044 => "0000000000000001000000000000100100000000000000111000101100011",
2045 => "0000000000000011000000000000001100000000000000111000101100101",
2046 => "0000000000000001000000000000000100000000000000011000101100111",
2047 => "0000000000000001000000000000001100000000000000111000101101010",
2048 => "0000000000000001000000000100101100000000000000111000101101101",
2049 => "0000000000000001000000000000001100000000000000011000101101111",
2050 => "0000000000000001000000000000001100000001000100101000101110001",
2051 => "0000000000000001000000000000001100000000000000111000101110011",
2052 => "0000000000000001000000000000001100000000000000111000101110101",
2053 => "0000000000000011000000000000001100000000000000011000101110111",
2054 => "0000000000000001000000000000010100000000000000111000101111001",
2055 => "0000001000100010000000000000001100000000000000011000101111011",
2056 => "0000000001000000000000000000001100000000001001011000101111101",
2057 => "0000000000000011000000000000001100000000000000111000101111111",
2058 => "0000000000000001000000000000001100000000000000011000110000001",
2059 => "0000000000000001000000000000001100000000010000011000110000011",
2060 => "0000000000000001000000010001000000000000000000111000110000101",
2061 => "0000000000000001000000000000001100000000000010011000110000111",
2062 => "0000000000010101000000000000100100000000000000111000110001010",
2063 => "0000000000000001000000000000100100000000000000111000110001100",
2064 => "0000000000000001000000000000001100000000000000011000110001110",
2065 => "0000000000000001000000000000001100000000000000111000110010000",
2066 => "0000000000000001000000000000000100000000000000111000110010010",
2067 => "0000000000000001000000000000100100000000000000111000110010100",
2068 => "0000000000000001000000000000001100000000000000011000110010111",
2069 => "0000000100010010000000000000010100000000000000111000110011001",
2070 => "0000010010001000000000000000000100000000000000111000110011011",
2071 => "0000000000000001000000000000101100000000000000111000110011110",
2072 => "0000000000000001000000000000000100000000000100111000110100000",
2073 => "0000000000000001000000000000000100000000000000111000110100011",
2074 => "0000000000000001000000000000010100000000000010011000110100110",
2075 => "0000000000000001000000000000001100000000001000111000110101001",
2076 => "0000000000000001000000001000101000000000000000111000110101011",
2077 => "0000000000000001000000000000000100000000000000111000110101110",
2078 => "0000000000000001000000000000001100000000000000111000110110000",
2079 => "0000000000000001000000000000001100000000101010111000110110010",
2080 => "0000000000000001000000000000001100000000101001001000110110100",
2081 => "0000000000000001000000000100001100000000000000111000110110110",
2082 => "0000000000000001000000000000000100000000000011111000110111000",
2083 => "0000000000000001000000000000001100000000000000011000110111010",
2084 => "0000000000000001000000000000001100000000100001001000110111100",
2085 => "0000000000000001000000000000001100000000000000111000110111111",
2086 => "0000000000000001000000000000001100000000000010011000111000001",
2087 => "0000000000000001000000000000001100000000010100001000111000011",
2088 => "0000000000000001000000000000000100000000000000011000111000101",
2089 => "0000000000000001000000000000001100000000010100111000111000111",
2090 => "0000000000000001000000000000001100000000100100001000111001010",
2091 => "0000000100101011000000000000001100000000000000111000111001101",
2092 => "0000000000000001000001010010100000000000000010111000111010000",
2093 => "0000000000000001000000000000001100000000000000111000111010011",
2094 => "0000000000000001000000000000100100000000000000111000111010101",
2095 => "0000000000010001000000000000001100000000000000111000111010111",
2096 => "0000000000000001000000000000000100000000000000111000111011010",
2097 => "0000000000000001000000000000010100000000000000111000111011101",
2098 => "0000000000000001000000000000001100000000000000011000111011111",
2099 => "0000000000010011000000000000001100000000000000011000111100001",
2100 => "0000000000000001000000000000001100000000000000011000111100011",
2101 => "0000000000100101000000000000001100000000000001011000111100101",
2102 => "0000000000000001000000010000000000000000000000111000111100111",
2103 => "0000000000000001000000010010100100000000000000111000111101010",
2104 => "0000000000000001000000000000000100000000000000111000111101101",
2105 => "0000000000000001000000000000001100000000000000111000111110000",
2106 => "0000000000000001000000000000101100000000001000111000111110011",
2107 => "0000000000000001000000000000001100000000000000011000111110110",
2108 => "0000000100100011000000000010001100000000000000111000111111000",
2109 => "0000000000000001000000000000001100000000100100001000111111010",
2110 => "0000000000000001000000000001010100000000000000111000111111100",
2111 => "0000000000000001000000000000010100000000000000111000111111110",
2112 => "0000000000000001000000000000001100000000000000011001000000000",
2113 => "0000000000000001000000000000010100000000000000111001000000010",
2114 => "0000000000000001000000001001001100000000000000111001000000100",
2115 => "0000000000000001000000000000001100000000000000111001000000110",
2116 => "0000000000000001000000000000000100000000000000011001000001000",
2117 => "0000000000000001000000000000001100000000000000111001000001010",
2118 => "0000000000000001000000000010010100000000000000111001000001100",
2119 => "0000000000000001000000000000001100000000000000111001000001110",
2120 => "0000000000000001000000000010100100000000000001011001000010000",
2121 => "0000000000000001000000000000001100000000000000011001000010010",
2122 => "0000000000000011000000000000001100000000000000011001000010100",
2123 => "0000000000000011000000000000001100000000000000111001000010110",
2124 => "0000010000010100000000000000001100000000100000111001000011000",
2125 => "0000000000000001000000000000001100000000000001011001000011010",
2126 => "0000000000000001000000000000000100000000000000111001000011100",
2127 => "0000000000000001000000000000001100000000000000111001000011110",
2128 => "0000000001000101000000000000000100000000000000111001000100000",
2129 => "0000000000000001000000000000001100000000000000111001000100010",
2130 => "0000000000000001000000000000001100000000000000011001000100100",
2131 => "0000000000000001000000000000001100000000000000011001000100110",
2132 => "0000000000000001000000000001001100000000000000111001000101000",
2133 => "0000000000000001000000000000001100000000000000011001000101010",
2134 => "0000000000000001000000000000101100000000000000111001000101100",
2135 => "0000000000000001000000000000001100000000000010111001000101110",
2136 => "0000000001000011000000000100100000000000000000111001000110000",
2137 => "0000000000000001000000000000000100000000000100001001000110010",
2138 => "0000000000000001000000000000001100000000000000011001000110100",
2139 => "0000000000000001000000000000000100000000000000111001000110110",
2140 => "0000000000000011000000000000000000000000000000111001000111000",
2141 => "0000000000000001000000000000000100000000000000111001000111010",
2142 => "0000000000000001000000000000001100000000000000111001000111100",
2143 => "0000000000000001000000000000001100000000000000011001000111111",
2144 => "0000000100100001000000000000001100000000000000111001001000001",
2145 => "0000000000000001000000000000001100000000000010101001001000011",
2146 => "0000000000000001000000000000000100000000000000111001001000101",
2147 => "0000000000000001000000000000000100000000000000111001001001000",
2148 => "0000000000001011000000000000001100000000000000111001001001010",
2149 => "0000000010100101000000000000001100000000100001011001001001100",
2150 => "0000000000000001000000000000001100000000000000011001001001110",
2151 => "0000000000000101000000000010101100000000000000111001001010000",
2152 => "0000000000000011000000000000000100000000000000111001001010010",
2153 => "0000000000000001000000000000000100000000000000111001001010100",
2154 => "0000000000000101000000000000000100000000000000111001001010111",
2155 => "0000000000000011000000000000001100000000000000111001001011001",
2156 => "0000000000000001000000000000001100000000000000111001001011011",
2157 => "0000000000000111000001000000000100000000001000101001001011101",
2158 => "0000000000000001000000000000001100000000000000111001001011111",
2159 => "0000000000001011000000000000000100000010101010101001001100001",
2160 => "0000000000000001000000000000001100000000000000111001001100011",
2161 => "0000000000000001000000000000001100000000000000011001001100101",
2162 => "0000000000000001000000000000001100000000000000011001001100111",
2163 => "0000000000000001000000010010100100000000000000011001001101001",
2164 => "0000000000000001000000000000001100000000000000111001001101011",
2165 => "0000000000000001000000000000001100000010000100011001001101110",
2166 => "0000000000000001000000000000000100000000000000111001001110001",
2167 => "0000000101010000000000000000001100000001010001011001001110100",
2168 => "0000000000000001000000000000001100000000000000111001001110111",
2169 => "0000000000000001000000000000000100000000000000111001001111001",
2170 => "0000000000000001000000010010010000000000000000111001001111011",
2171 => "0000000000000001000000000000001100000000000000011001001111110",
2172 => "0000000000000001000000000000001100000000000000111001010000000",
2173 => "0000000000000001000000000000100100000000000000011001010000010",
2174 => "0000000000000001000000000000001100000000000000011001010000100",
2175 => "0000000000000001000000000000000100000000000000111001010000111",
2176 => "0000000000000001000000000000000100000000000000111001010001001",
2177 => "0000000010100001000000000001010000000000000000011001010001011",
2178 => "0000000000000001000000000000001100000000000000111001010001101",
2179 => "0000000000000001000000000000010100000000000000111001010001111",
2180 => "0000010100100101000000000000001100000000010010111001010010001",
2181 => "0000001000010000000000000000000000000000000000011001010010011",
2182 => "0000000000000001000000000101000100000000000000111001010010110",
2183 => "0000000000000001000000000001010100000000000010101001010011000",
2184 => "0000000000000001000000000000001100000000000000111001010011010",
2185 => "0000000000000001000000000000001100000000000101011001010011100",
2186 => "0000000001000001000000000000001100000000001000111001010011110",
2187 => "0000000000000001000000001000010100000000000000111001010100001",
2188 => "0000000000000001000000000000001100000000000000011001010100011",
2189 => "0000000010010001000000000000001100000000000000111001010100101",
2190 => "0100010000000100000000000000001100000000000000011001010101000",
2191 => "0000000000000001000000000000001100000000000000011001010101010",
2192 => "0000000000000001000000000000001100000000000000011001010101100",
2193 => "0000000000000001000000000010101000000000000100111001010101111",
2194 => "0000000000000001000000000000000100000000000000111001010110001",
2195 => "0000000000000001000000000000100100000000000000111001010110011",
2196 => "0000000000000101000000000000001100000000100000011001010110101",
2197 => "0000000000000001000000000000101100000000000100101001010110111",
2198 => "0000000000000001000000001001001100000000000000111001010111010",
2199 => "0000000000000001000000000010100100000000000000111001010111100",
2200 => "0000000000000001000000000101000000000000000000111001010111111",
2201 => "0000000000000001000000000000001100000000000000111001011000001",
2202 => "0000000000000001000000000000001100000000000000111001011000011",
2203 => "0000000000001001000000000000000100000000000000111001011000101",
2204 => "0000000000000001000000000000000100000000000000111001011000111",
2205 => "0000000000000011000000000000000100000000000000111001011001010",
2206 => "0000001000001001000000000000001100000000000000111001011001101",
2207 => "0000000000000001000000000000001100000000000000011001011010000",
2208 => "0000000100100011000000000000001100000000000000111001011010010",
2209 => "0000000000000001000000000010000100000000000000111001011010100",
2210 => "0000000000000001000000000000000100000000000000111001011010110",
2211 => "0000000000000001000000001010010100000000000000111001011011000",
2212 => "0000000000000001000000000000010100000000000000111001011011010",
2213 => "0000000000000001000000000000001100000000000100111001011011100",
2214 => "0000000000000001000000000000001100000000000000111001011011110",
2215 => "0000000000000001000000000000001100000001010100001001011100000",
2216 => "0000000000000001000000000000001100000000000000111001011100010",
2217 => "0000000000000001000000000000001100000000000000111001011100100",
2218 => "0000000000001011000000000000001100000000000010011001011100110",
2219 => "0000000000000011000000000000000100000000000000111001011101000",
2220 => "0000000000000001000000000000000100000000000000111001011101010",
2221 => "0000000000000001000000000000001100000000000000011001011101100",
2222 => "0000000000000001000000000000001100000000000001011001011101110",
2223 => "0000000100100101000000000000001100000000000000111001011110000",
2224 => "0000000000000001000000000000001100000000000000111001011110010",
2225 => "0000000001010101000000000000001100000000000000111001011110100",
2226 => "0000000000000001000000000000001100000000000010011001011110110",
2227 => "0000000000000001000000000000000100000000000000011001011111000",
2228 => "0000000000000001000000000000010100000000000000111001011111010",
2229 => "0000000000000011000000000000100100000000000000111001011111100",
2230 => "0000000000000001000000000000001100000000000000011001011111110",
2231 => "0000000000000001000000000000001100000000001010111001100000001",
2232 => "0000000000000001000000000000001100000000000000111001100000011",
2233 => "0000000000000001000000000000000100000000000100011001100000101",
2234 => "0000000000000001000000000000000100000000000000111001100000111",
2235 => "0000000000000001000000000000000100000000010000101001100001001",
2236 => "0000000000000001000000000000001100000001000001011001100001011",
2237 => "0000000000000001000000001010100000000000000000111001100001101",
2238 => "0000000000000001000000000000001100000000000000011001100001111",
2239 => "0000000000011011000000000000001100000000000000011001100010010",
2240 => "0000000000000001000000000000001100000000000000111001100010100",
2241 => "0000000000000001000000000000001100000000000000111001100010110",
2242 => "0000000000000101000000000000001100000000000000111001100011000",
2243 => "0000000000000001000000000000001100000000001001011001100011010",
2244 => "0000000100000011000000000000001100000000000000011001100011100",
2245 => "0000010010101000000000000100100100000000000000111001100011110",
2246 => "0000000000100001000000000000001100000000000000011001100100001",
2247 => "0000000000000001000000000000000100000000010000101001100100011",
2248 => "0000000000000001000000000000000100000000000000111001100100101",
2249 => "0000000000000001000000000000001100000000000100011001100100111",
2250 => "0000000000000001000000000000000100000000000000111001100101001",
2251 => "0000000000000101000000000000001100000000000000011001100101011",
2252 => "0000000000000011000000000000010100000000000000111001100101101",
2253 => "0000000000000001000000000000000100000000000001011001100110000",
2254 => "0000000000000011000000000000001100001001001010001001100110011",
2255 => "0000000000000001000000000000000100000000000000111001100110101",
2256 => "0000000000000001000000000000001100000000000000111001100110111",
2257 => "0000000000000001000001010010010000000000000000011001100111001",
2258 => "0000000000000001000000000000001100000000000000111001100111011",
2259 => "0000000000000001000000000000000100000000000000111001100111101",
2260 => "0000001000001001000000000000001100000000000000111001100111111",
2261 => "0000010010000001000000000000101100000000000000111001101000001",
2262 => "0000000000000001000000000000001100000000000000111001101000011",
2263 => "0001000010000011000000000100001100000000000000111001101000101",
2264 => "0000000000000001000000000000001100000000000000111001101000111",
2265 => "0000000000000001000000000000000100000000000000111001101001010",
2266 => "0000000000000001000000000000001100000000000010111001101001101",
2267 => "0000000000000001000000000000001100000000101001001001101001111",
2268 => "0000000100010100000000000000001100000010010000011001101010001",
2269 => "0000000000000001000000000000001100000000000000011001101010011",
2270 => "0000000000000011000000000000001100000000000000011001101010101",
2271 => "0000000001000001000000001010010100000000000000111001101010111",
2272 => "0000000000000001000000000000001100000001000001011001101011001",
2273 => "0000000000000001000000000000000100000000001000001001101011011",
2274 => "0000000000000001000000000000001100000000000000111001101011110",
2275 => "0000000000000001000000000000000100000000000000111001101100000",
2276 => "0000000000000001000000000000001100000000000000111001101100011",
2277 => "0000000000000001000000001000010000000000000000111001101100101",
2278 => "0000000000000001000000000000001100000000000000111001101100111",
2279 => "0000000000000001000000000000000100000000000000111001101101010",
2280 => "0000000000000001000000000000000100000000000000111001101101101",
2281 => "0000000000000001000000000000001100000000001001011001101101111",
2282 => "0000000000000001000000000000001100000000000000111001101110001",
2283 => "0000000000000101000000001000100100000000000000111001101110011",
2284 => "0000000000000111000000001000001100000000000000111001101110101",
2285 => "0000000000000101000000000000001100000000000000011001101110111",
2286 => "0000000000000001000000000000000100000000000000111001101111001",
2287 => "0000000000000001000000000000010100000000000000011001101111011",
2288 => "0000000000000101000000000000001100000000000000011001101111110",
2289 => "0000000000000001000000000000000100000000000000111001110000000",
2290 => "0000000000010101000000000000001100000000000000011001110000011",
2291 => "0000000000000001000000000000001100000000000001011001110000110",
2292 => "0000000000000001000000000000001100000000000000011001110001001",
2293 => "0000000000000001000000000000010100000000000000111001110001100",
2294 => "0000000000100101000000000000001100000000000000111001110001110",
2295 => "0000000000000001000000000000001100000000000000011001110010000",
2296 => "0000000000001011000000000000001100000000000000111001110010010",
2297 => "0000001000001010000000000001010100000000000000111001110010100",
2298 => "0000010001010100000000000000001100000001001001011001110010110",
2299 => "0000000000000001000000001001010100000000000000011001110011000",
2300 => "0000000000001001000000000000001100000000000000011001110011010",
2301 => "0000000000000001000000000000000100000000000000011001110011100",
2302 => "0000000000000001000000000000000100000000000000111001110011110",
2303 => "0000000000000011000000000000001100000000000100111001110100000",
2304 => "0000000000000001000000000000001100000000000001011001110100010",
2305 => "0000000000000001000000000000001100000000000000011001110100100",
2306 => "0000000000000001000000000000001100000000000100111001110100110",
2307 => "0000000000000101000000000000001100000000001010011001110101000",
2308 => "0000000000000001000000000000001100000000000000111001110101010",
2309 => "0000000000000001000000000000000100000000000000111001110101100",
2310 => "0000000000000001000000000000001100000000000100011001110101110",
2311 => "0000000000001011000000000010100000000000000000111001110110000",
2312 => "0000001010000010000000000000001100000000000000011001110110010",
2313 => "0000000000000001000000000000001100000000000000111001110110100",
2314 => "0000000000000001000000000010101100000000000000111001110110110",
2315 => "0000000000100011000000000000001100000000000000011001110111000",
2316 => "0000000000100101000000000000000100000000000000111001110111010",
2317 => "0000000000000001000000000000010100000000000000111001110111100",
2318 => "0000000000000001000000000000001100000000100001001001110111110",
2319 => "0000000000000001000000000000001100000000000000011001111000001",
2320 => "0000000000000101000000000100010100000000000000111001111000011",
2321 => "0000000000000001000000000000001100000000000000111001111000110",
2322 => "0000000000000001000000000000001100000000100010011001111001001",
2323 => "0000000000001001000000000000001100000000000000011001111001100",
2324 => "0000000000000001000000000000010100000000000000111001111001110",
2325 => "0000000000000001000000000000001100000000000000111001111010000",
2326 => "0000000010010010000000000000001100000000000000011001111010010",
2327 => "0000000000000001000000000000001100000000000000111001111010100",
2328 => "0000000000000001000000000000001100000000001000011001111010110",
2329 => "0000001001010100000000000000001100000000001000011001111011000",
2330 => "0000000000000001000000000000001100000000000001011001111011011",
2331 => "0000000000000001000000000000001100000000000000101001111011101",
2332 => "0000000000001001000000000000000100000000000000111001111011111",
2333 => "0000000000000001000001000010000000000000000000111001111100001",
2334 => "0000000000000001000000000000000100000000001010001001111100011",
2335 => "0000000000000001000000000000001100000000000000111001111100101",
2336 => "0000000000000001000000100101000000000000000000111001111100111",
2337 => "0000000000000001000000000000001100000000000010011001111101001",
2338 => "0000000000000001000000000000001100000000000000011001111101100",
2339 => "0000000000000101000000000000001100000000000000111001111101111",
2340 => "0000000000000001000000000000000100000000000000111001111110010",
2341 => "0000000000000001000000000010101100000000000000111001111110100",
2342 => "0000000000000011000000000000001100000000000000111001111110111",
2343 => "0000000000000001000000000000001100000000000000111001111111001",
2344 => "0000000000000001000000000000001100000000000100111001111111011",
2345 => "0000000000000001000000000000000100000000000000111001111111101",
2346 => "0000000000000001000000000000100100000000000000111001111111111",
2347 => "0000000000000001000000000000001100000000001000111010000000010",
2348 => "0000000000000001000000000000001100000000000010111010000000101",
2349 => "0000000000000001000000000000001100000000100000011010000000111",
2350 => "0000000000000001000000000000000100000000000000111010000001001",
2351 => "0000000000001001000000000000100100000000000000111010000001100",
2352 => "0000000000001001000000000000000100000000001000111010000001111",
2353 => "0000000100001011000000000000001100000000000000011010000010001",
2354 => "0000000000000001000000000000000100000000000100011010000010011",
2355 => "0000000000000001000000000000010100000000000000111010000010110",
2356 => "0000000000000001000000000000001100000000000010111010000011000",
2357 => "0000000000000001000000100001000000000000000000111010000011011",
2358 => "0000000000010001000000000000100100000000000000111010000011101",
2359 => "0000000000000001000000000000001100000000000000111010000011111",
2360 => "0000000000000001000000000000000100000000000000111010000100001",
2361 => "0000000000000001000000000000000100000000000000111010000100011",
2362 => "0000000000000001000000000000001100000000000000111010000100101",
2363 => "0000000000000001000000000000000100000000000000111010000100111",
2364 => "0000000000000001000000000000010100000000000000011010000101001",
2365 => "0000000000000001000000000000000100000000000000111010000101011",
2366 => "0000000000000001000000000000001100000000000000011010000101110",
2367 => "0000000000000001000000000000001100000000000000011010000110000",
2368 => "0000000000000001000000000000000100000000000000011010000110010",
2369 => "0000000000000001000000000000000100000000000000111010000110101",
2370 => "0000000000000001000000000000000100000000000000111010000111000",
2371 => "0000000000000001000000000001001100000000000000111010000111010",
2372 => "0000000000000001000000000000001100000000000101011010000111100",
2373 => "0000000000000001000000000000001100000000000000111010000111110",
2374 => "0000000000000001000000000000000100000000000000111010001000000",
2375 => "0000000000000001000000000000001100000000000000111010001000011",
2376 => "0000000000000001000000000000001100000000000000111010001000101",
2377 => "0000000000000001000000000000001100000000000001011010001000111",
2378 => "0000000000000001000000000000001100000000000000011010001001001",
2379 => "0000000000000001000000000010010100000000000000111010001001100",
2380 => "0000000101010010000000000000001100000000000000011010001001110",
2381 => "0000000000000001000000000000000100000000000000111010001010000",
2382 => "0000010010100101000000000000000110001000000000001010001010010",
2383 => "0000000000000001000000000000001100000000000000111010001010101",
2384 => "0000000000000001000000001000101000000000000000111010001011000",
2385 => "0000000000000101000000000000001100000000000000011010001011010",
2386 => "0000000000000001000000000000001100000000000000011010001011100",
2387 => "0000000000000001000000000000000100000000000000111010001011111",
2388 => "0000000000000001000000000000000100000000000000001010001100001",
2389 => "0000000000000001000000000000001100000000000000111010001100011",
2390 => "0000000000100001000000000010010100000000000000111010001100101",
2391 => "0000000000000001000000000100000100000000000000111010001100111",
2392 => "0000000000000001000000000000001100000000000000111010001101001",
2393 => "0000000000000001000000000000001100000000000000011010001101011",
2394 => "0000000000000001000000000000001100000000000001011010001101101",
2395 => "0000000000000001000000010000000100000000000000111010001101111",
2396 => "0000000000000001000000000000000100000000010010101010001110010",
2397 => "0000000000001001000000000000001100000000000000111010001110100",
2398 => "0000000000000001000000000000001100000000000000111010001110110",
2399 => "0000000000000011000000000100010000000000000000111010001111000",
2400 => "0000010010000101000000001001001000000000000000111010001111010",
2401 => "0000000000000001000000000000001100000000000000111010001111100",
2402 => "0000000000000001000000000000001100000001001001011010001111110",
2403 => "0000000000000001000000000000001100000000000000111010010000000",
2404 => "0000010101001001000000000001000100000000000000111010010000010",
2405 => "0000000000000001000000000000001100000000000000111010010000100",
2406 => "0000000000000001000000000000010100000000000000111010010000110",
2407 => "0000000000000001000000000000001100000000000000111010010001000",
2408 => "0000000000000001000000000000100100000000010101011010010001010",
2409 => "0000000000000001000000000000000100000000000000111010010001100",
2410 => "0000000000000001000000000000001100000000010000011010010001110",
2411 => "0000000000000001000000000000000100000000000000111010010010000",
2412 => "0000000000000001000000000000001100000000000000011010010010010",
2413 => "0000000000000001000000000000001100000000000000111010010010101",
2414 => "0000000000001001000000000000000100000000000000011010010010111",
2415 => "0000000000000001000000000000001100000000000000011010010011001",
2416 => "0000000000000001000000000000001100000000100010001010010011011",
2417 => "0000000000000001000000000000001100000010010101011010010011101",
2418 => "0000001001010001000000001000100000000000000000111010010011111",
2419 => "0000000000000001000000000000001100000000000000111010010100001",
2420 => "0000000000000011000000000000000100000000000001011010010100011",
2421 => "0000000000000001000000001010001000000000000000111010010100101",
2422 => "0000000000000001000000000000001100000000000000011010010100111",
2423 => "0000000000000001000000000000001100000000000000011010010101001",
2424 => "0000000000000001000000000000001100000000000000011010010101011",
2425 => "0000000000000001000000000000001100000000000101001010010101101",
2426 => "0000000000000001000000000000001100000000000100011010010110000",
2427 => "0000000000000001000000001000010100000000000000111010010110010",
2428 => "0000000000000001000000000000001100000000010100011010010110100",
2429 => "0000000000000001000000000000000100000000000000111010010110111",
2430 => "0000000000000001000000000000000100000000000000111010010111010",
2431 => "0000000000000101000000000000001100000000000000111010010111100",
2432 => "0000000000000001000000000000000100000000000000111010010111110",
2433 => "0000000000000001000000000000001100000000000000111010011000000",
2434 => "0000000000000001000000000000001100000000000000011010011000011",
2435 => "0000000000010101000000000000001100000000000000111010011000101",
2436 => "0000000000000001000000000000000100000000000000111010011000111",
2437 => "0000001000100000000000000000001100000100100010001010011001010",
2438 => "0000000000000101000000000000101100000000000000011010011001101",
2439 => "0000000000000001000000000000001100000000000000111010011010000",
2440 => "0000000000000001000000000001001100000000000000111010011010010",
2441 => "0000000000000001000000000000001100000000001010111010011010100",
2442 => "0000000000000101000000000000010100000000000000111010011010111",
2443 => "0000000000000001000000000000000100000000000000111010011011001",
2444 => "0000000000000001000000000000001100000000001001011010011011011",
2445 => "0000000000010011000000000000001100000000000000111010011011101",
2446 => "0000000000000001000000000000000100000000000000011010011100000",
2447 => "0000000000000001000000000000000100000000000000111010011100010",
2448 => "0000000000000001000000000000001100000000000000011010011100100",
2449 => "0000000000101011000000000000001100000001000001011010011100111",
2450 => "0000000000000001000000000000010100000000010010001010011101001",
2451 => "0000000000000001000000000000001100000000101000001010011101011",
2452 => "0000000000000001000000000000100100000000000000111010011101101",
2453 => "0000000000000001000000000000001100000000000000011010011101111",
2454 => "0000000000000001000000000000000100000000000000111010011110001",
2455 => "0000000000000001000000000000000100000000000000111010011110011",
2456 => "0000000000000001000000001000010000000000000000111010011110101",
2457 => "0000000000000101000000000000001100000000000000111010011111000",
2458 => "0000000000000001000000000000001100000000010100011010011111011",
2459 => "0000000000000101000000000000010000000000000000111010011111101",
2460 => "0000000000000001000000000001010100000000000000111010011111111",
2461 => "0000000000000001000000100101001100000000000000111010100000010",
2462 => "0000000000000001000000000000001100000000000000111010100000100",
2463 => "0000000100101001000000000000001100000000000001011010100000110",
2464 => "0000000000000001000000000000000000000000000000011010100001001",
2465 => "0000000000000001000000000000001100000101000000101010100001011",
2466 => "0000000000000001000000000000001100000000100100011010100001101",
2467 => "0000000000000011000000000000001100000000000001011010100001111",
2468 => "0000010100010011000000000100101100000000000000111010100010001",
2469 => "0000000000010001000000000000001100000000000000111010100010011",
2470 => "0000000000000001000000000000101100000000000000011010100010101",
2471 => "0000000000000001000000000000010100000000000000111010100010111",
2472 => "0000000000000001000000000000001100000001010001001010100011001",
2473 => "0000000000000001000000000000001100000000000101011010100011011",
2474 => "0000000000000001000000000000001100000000000000011010100011101",
2475 => "0000000000000001000000000000001100000000000101001010100011111",
2476 => "0000000000000001000000000000000100000000001000101010100100001",
2477 => "0000000000000001000000000001000100000000000000111010100100011",
2478 => "0000000000000001000000000010010100000000000000011010100100101",
2479 => "0000000000000001000000000000001100000000000001011010100100111",
2480 => "0000000000000101000000000000010100000000000000111010100101010",
2481 => "0000000000100101000000000000001100000000000010111010100101100",
2482 => "0000000101000000000000000000000100000000000000011010100101110",
2483 => "0000000000000001000000000000001100000000000000111010100110000",
2484 => "0000000000000001000000000000001100000000010000101010100110010",
2485 => "0000000000000001000000000000010100000000000000111010100110100",
2486 => "0000000000000001000000000000001100000000100000101010100110111",
2487 => "0000000000000001000000000000001100000000000000111010100111001",
2488 => "0000000000000001100010000000000000000000000000011010100111011",
2489 => "0000000000000001000000000000001100000000000000111010100111101",
2490 => "0000000000000011000000000000001100000000000010011010100111111",
2491 => "0000000000000001000000000000001100000100010100101010101000010",
2492 => "0000000000010001000000000000001100000000000000011010101000101",
2493 => "0000000000000001000000000000001100000000000000011010101001000",
2494 => "0000000000000001000000000010001100000000000000011010101001011",
2495 => "0000000010100010000000000000001100000000000000011010101001101",
2496 => "0000000000000001000000000000100100000000000000111010101001111",
2497 => "0000000000000001000000000000001100000000000100011010101010010",
2498 => "0000000000001001000000000001001100000000000000111010101010100",
2499 => "0000000010100001000000000000000100000000000000111010101010110",
2500 => "0000000000000001000000000101000100000000010000011010101011000",
2501 => "0000000000000001000000000000001100000000000000011010101011010",
2502 => "0000000000101011000000000000001100000000000000011010101011101",
2503 => "0000000000001001000000000000001100000000000000011010101011111",
2504 => "0000000000101001000000000000001100000000000000011010101100001",
2505 => "0000000000000001000000000010000100000000000000111010101100011",
2506 => "0000000000000101000000000000001100000000000010011010101100101",
2507 => "0000000000000001000000000000001100000000000000011010101100111",
2508 => "0000000000000001000000000000000100000000000000111010101101001",
2509 => "0000000000000101000000000000001100000000000000111010101101011",
2510 => "0000000000000001000000000000001100000000000010011010101101101",
2511 => "0000000000000001000000000000000100000000000000111010101110000",
2512 => "0000000000000001000000000010101100000000000000111010101110011",
2513 => "0000000000000011000000000000000100000000000000111010101110101",
2514 => "0000000000010011000000000000001100000000000000111010101111000",
2515 => "0000000000000001000000000000100100000000000000111010101111010",
2516 => "0000000000000101000000000000000100000000000000111010101111100",
2517 => "0000000000000001000000000000001100000000000000011010101111110",
2518 => "0000000000000001000000000000001100000000000000111010110000000",
2519 => "0000000000000001000000000000010100000000000000111010110000010",
2520 => "0000000000000001000000000000001100000000000000111010110000100",
2521 => "0000000000000001000000000000001100000000000001011010110000110",
2522 => "0000000000000001000000000000000100000000000000111010110001000",
2523 => "0000000000000001000000000000001100000000000001011010110001010",
2524 => "0000000000000001000000000000001100000000000000111010110001100",
2525 => "0000000000000001000000001010101000000000000000111010110001110",
2526 => "0000000000000001000000000000001100000000000000111010110010000",
2527 => "0000000000000001000000000001000100000000000000111010110010010",
2528 => "0000000000000001000000000010010100000000000000111010110010100",
2529 => "0000000000000001000000000000001100000000000000011010110010110",
2530 => "0000000000000001000000001001001100000000000000111010110011000",
2531 => "0000000000000001000000000000001100000000001000011010110011010",
2532 => "0000001010100010000000000000001100000010001010001010110011100",
2533 => "0000000000000001000000000000101100000000000000111010110011110",
2534 => "0000000000000001000000000000001100000000000000011010110100000",
2535 => "0000000000000001000000000010100100000000000000111010110100010",
2536 => "0000000000000001000000000001000100000000000000111010110100101",
2537 => "0000000000000001000000001000000100000000000000111010110101000",
2538 => "0000000000000001000000000000000100000000000000111010110101011",
2539 => "0000000000000001000000000000001100000000000000111010110101101",
2540 => "0000000000000001000000000000101100000000000000111010110110000",
2541 => "0000000000000001000000000000001100000000000000011010110110011",
2542 => "0000000000000001000000000000001100000000001000011010110110101",
2543 => "0000000000000001000001010010010000000000000001011010110111000",
2544 => "0000000000000001000000000000000100000000000000111010110111011",
2545 => "0000000000010001000000000000000110001000000000001010110111110",
2546 => "0000000000000001000000000000001100000000000000111010111000000",
2547 => "0000000000000001000000000000001100000000101000001010111000010",
2548 => "0000000000000001000000000000000100000000000000111010111000100",
2549 => "0000000000000001000000000000001100000000000000111010111000110",
2550 => "0000000000000001000000000001001100000000000000111010111001000",
2551 => "0000000000010101000000000000001100000000000000011010111001010",
2552 => "0000000000000001000000000000000100000000000000111010111001100",
2553 => "0000000000000001000000000000001100000010100101011010111001110",
2554 => "0000000000000001000000000000001100000000000000111010111010001",
2555 => "0000000000000001000000000000001100000000000000011010111010011",
2556 => "0000000000000001000000000000000100000000000000111010111010110",
2557 => "0000000000000001000000000000001100000000000001011010111011000",
2558 => "0000000000000001000000000000001100000010000000011010111011010",
2559 => "0000000000000001000000000000000100000000000000111010111011100",
2560 => "0000000000000001000000010000000000000000000000111010111011110",
2561 => "0000000000000001000000000001000100000000000000111010111100000",
2562 => "0000000000000001000000000000001100000000000000111010111100010",
2563 => "0000000000000001000000000001001100000000010101001010111100100",
2564 => "0000000000000001000000000000000100000000000000111010111100110",
2565 => "0000000000000001000000000001001100000000000000111010111101000",
2566 => "0000000000000001000000000000001100000000000000111010111101010",
2567 => "0000000101010001000000000000001100000000000000111010111101100",
2568 => "0000000000000001000000000000001100000000000000111010111101110",
2569 => "0000000000000101000000000000001100000000000101011010111110001",
2570 => "0000000000000001000000000000001100000000000100111010111110011",
2571 => "0000000000000011000000000010010100000000000000111010111110101",
2572 => "0000000000000001000000000000001100000000000000111010111110111",
2573 => "0000000010000001000000000000000100000000000000111010111111001",
2574 => "0000000000000001000000000000001100000000000000111010111111011",
2575 => "0000000000000001000000000000001100000000000001011010111111101",
2576 => "0000000000000001000000000000001100000000000000111010111111111",
2577 => "0000000000000001000000000000001100000000000000011011000000001",
2578 => "0000000000000001000000000000100100000000000000111011000000011",
2579 => "0000000000000011000000000000010000000000000000111011000000101",
2580 => "0000000000000001000000000000001100000000001000011011000000111",
2581 => "0000000000000001000000000101001100000000000000111011000001010",
2582 => "0000000000000101000000000000001100000000000001011011000001101",
2583 => "0000000000000001000000000000001100000000000000111011000010000",
2584 => "0000000000000001000000000000001100000000000000111011000010011",
2585 => "0000000000000001000000000000001100000000000001011011000010110",
2586 => "0000000000000101000000000000001100000000000000011011000011000",
2587 => "0000000000000001000000000000001100000000000000011011000011010",
2588 => "0000000000000001000000001000101100000000000000111011000011101",
2589 => "0000000000000001000000000000000100000000000000111011000011111",
2590 => "0000000000000001000000010000100100000000000000111011000100010",
2591 => "0000000000000001000000000000001100000000000000011011000100101",
2592 => "0000000000001011000000000000100100000000000000111011000100111",
2593 => "0000010000010101000000000000000100000000000000111011000101010",
2594 => "0000000000000001000000000000101100000000000000111011000101100",
2595 => "0000000000000001000000010101000100000000000000111011000101110",
2596 => "0000000000000001000000000000001100000000000100011011000110001",
2597 => "0000000000000001000000000000100100000000000000111011000110011",
2598 => "0000000000000001000000000000001100000000000000111011000110110",
2599 => "0000000000000001000000000000000100000000000000111011000111001",
2600 => "0000000000000001000000000000001100000000000000111011000111011",
2601 => "0000000010000100000000000000001100000000001000011011000111101",
2602 => "0000000000000001000000000000001100000000000000011011000111111",
2603 => "0000000000000001000000101010101000000000000000011011001000001",
2604 => "0000000000001001000000000000001100000000000010011011001000011",
2605 => "0000000000000011000000001000010100000000000000111011001000101",
2606 => "0000000000000001000000000000001100000000000000111011001000111",
2607 => "0000000000000001000000000000001100000000000000111011001001001",
2608 => "0000000000000001000000000000000100000000000000111011001001011",
2609 => "0000000000001001000000000000001100000000000000111011001001110",
2610 => "0000000000000001000000000000001100000000000000111011001010000",
2611 => "0000000000000001000000000000100100000000000000111011001010010",
2612 => "0000100001000001000000000000001100001010001010101011001010101",
2613 => "0000000000000001000000000000001100000000001001011011001011000",
2614 => "0000000000000011000000000000001100000000000101011011001011010",
2615 => "0000000000000001000000000000001100000001000101001011001011100",
2616 => "0000000000000001000000010010101000000000000000111011001011110",
2617 => "0000000000000001000000000000000100000000000000011011001100001",
2618 => "0000000000000001000000000000001100000000000000011011001100011",
2619 => "0000000000000001000000000000001100000000001000011011001100101",
2620 => "0000000000000001000000000000001100000000010010001011001100111",
2621 => "0000000000000001000000000000001100000000000010111011001101001",
2622 => "0000000000000001000000000000000100000000000000111011001101011",
2623 => "0000000000000101000000000000000100000000000001011011001101101",
2624 => "0000000000000011000000000000001100000000000001011011001101111",
2625 => "0000000000000001000000010000000000000000000000111011001110001",
2626 => "0000000000000101000000000000001100000000000000011011001110011",
2627 => "0000000000000101000000000001010100000000000000111011001110110",
2628 => "0000001010010001000000000000001100000000000000111011001111000",
2629 => "0000000000000001000000000000001100000000000000011011001111010",
2630 => "0000000000000001000000000000001100000000000000011011001111100",
2631 => "0000000000000001000000000001000100000000010000111011001111110",
2632 => "0000000000000001000000000000001100000000001000111011010000000",
2633 => "0000000000000001000000000000001100000000000000011011010000010",
2634 => "0000000000000001000000000000001100000000000000111011010000100",
2635 => "0000000000000011000000000100001100000000000000111011010000110",
2636 => "0000000000000001000000000000001100000000000000111011010001000",
2637 => "0000000001010001000000000000000100000000000010011011010001010",
2638 => "0000000000000011000000000000001100000000000000011011010001100",
2639 => "0000000000000001000000000000001100000000000000011011010001110",
2640 => "0000000000000001000000000000010100000000000000111011010010000",
2641 => "0000000000000001000000000000000100000000000000111011010010010",
2642 => "0000000010000010000000000000001100000000000101011011010010101",
2643 => "0000000000000001000000000000001100000000000101011011010011000",
2644 => "0000000000000001000000000000000100000000000000111011010011010",
2645 => "0000000000000001000000000000001100000000100000101011010011100",
2646 => "0000000000001001000000000000001100000000000000111011010011111",
2647 => "0000000000001011000000000000000100000000000011111011010100010",
2648 => "0000000000000001000000000000001100000000000000111011010100100",
2649 => "0000000000010101000000000000001100000000000001011011010100111",
2650 => "0000000000010011000000000010100100000000000000111011010101001",
2651 => "0000000000000001000000000000001100000000000000011011010101011",
2652 => "0000100101000010000000000000001100000000000000111011010101101",
2653 => "0000000000000001000000000000000100000000000010111011010101111",
2654 => "0000000000000001000000000000001100000000001010111011010110010",
2655 => "0000000000000001000000000010010100000000000000111011010110100",
2656 => "0000000000000001000000000000001100000000000000011011010110110",
2657 => "0000000000000001000000000000001100000000000000111011010111001",
2658 => "0000000000000001000000000000001100000000000000011011010111011",
2659 => "0000000000000001000000000000000100000000000000111011010111101",
2660 => "0000000000000001000000000000001100000000000000111011010111111",
2661 => "0000000000000100000000000000001100000000000000011011011000001",
2662 => "0000000000000001000000001010100100000000000000111011011000011",
2663 => "0000000000000001000000000000001100000000010001011011011000101",
2664 => "0000000000000001000000000000001100000000000000011011011000111",
2665 => "0000000000000011000000000000000100000000000000111011011001001",
2666 => "0000000000000001000000000000000100000000000000111011011001011",
2667 => "0000101001000000000000000000000100000000000000111011011001101",
2668 => "0000000001010001000000000000001100000000000101011011011001111",
2669 => "0000000101010011000000000000000100000000000000111011011010001",
2670 => "0000000000000001000000000001010100000000000000111011011010011",
2671 => "0000000000000011000000001010001000000000000000111011011010110",
2672 => "0000101000001010000000000000001100000000000000111011011011001",
2673 => "0000000000010001000000000000000100000000000000111011011011011",
2674 => "0000000000000001000000000000001100000000000000111011011011101",
2675 => "0000000000001001000000000000000100000000000000111011011100000",
2676 => "0000000101001001000000000000001100000000000000011011011100011",
2677 => "0000000000010001000000000000000100000000000000111011011100101",
2678 => "0000000000000001000000000000001100000000000000111011011100111",
2679 => "0000000000000001000000000000001100000000000000111011011101001",
2680 => "0000000000000001000000000000001100000000000000011011011101100",
2681 => "0000000000000001000000000000000100000000000000111011011101110",
2682 => "0000000010100101000000000000001100000000000000111011011110000",
2683 => "0000000000000001000000000000001100000000101001001011011110010",
2684 => "0000000000000001000000000000001100000000000001001011011110100",
2685 => "0000000000000001000000000000001100000000001000111011011110110",
2686 => "0000000000000001000000000000000100000000000000111011011111000",
2687 => "0000000000000101000000000000000100000000000010011011011111010",
2688 => "0000000000010101000000000000001100000000000000111011011111100",
2689 => "0000000000000001000000000100100000000000010010111011011111110",
2690 => "0000000000000011000000000000001100000000000000011011100000000",
2691 => "0000000000000001111010100100000000000000000000011011100000010",
2692 => "0000000000000001000000000000000100000000000000111011100000100",
2693 => "0000000000010101000000000000001100000000000000111011100000110",
2694 => "0000000000000001000000000000001100000000000000011011100001000",
2695 => "0000000000000001000000000000000100000000000001011011100001010",
2696 => "0000000000000001000000000000001100000000000000111011100001100",
2697 => "0000000000001011000000000000001100000000000000011011100001110",
2698 => "0000000000000001000000000000001100000000000000111011100010000",
2699 => "0000001000001001000000000000000100000000000000111011100010010",
2700 => "0000101010010001000000000000001100000000000000111011100010100",
2701 => "0000000000001011000000000001000100000001010010001011100010110",
2702 => "0000000000000001000000000000001100000000000000011011100011000",
2703 => "0000000001001011000000000000001100000000000010011011100011010",
2704 => "0000000000000001000000000000001100000000010001011011100011100",
2705 => "0000000000000001000000001000000100000000000000111011100011110",
2706 => "0000000000000001000000000000001100000000000000111011100100000",
2707 => "0000000000000001000000000000001100000000000000011011100100011",
2708 => "0000000000000001000000000000001100000000000000111011100100110",
2709 => "0000000000000001000000000000001100000000000010111011100101000",
2710 => "0000000000000001000000000000001100000000000000111011100101010",
2711 => "0000000000000001000000000000010100000010100100011011100101100",
2712 => "0000000000000001000000000000000100000000000000111011100101111",
2713 => "0000000000000001000000000000010100000000000000111011100110001",
2714 => "0000000001000101000000000000001100000000000000011011100110011",
2715 => "0000000000000001000000000000001100000000000000011011100110101",
2716 => "0000000000000011000000000000000100000000000000111011100110111",
2717 => "0000000000000001000000000000001100000000000000111011100111001",
2718 => "0000000000000101000000000000001100000000000000011011100111011",
2719 => "0000000000000001000000000000101100000000000000111011100111110",
2720 => "0000000000000001000000000000001100000000000101011011101000000",
2721 => "0000000000000001000000000001000100000000000000111011101000010",
2722 => "0000000000000001000000000000001100000001000001001011101000100",
2723 => "0000001000010100000000000000010100000000000000111011101000110",
2724 => "0000000000000101000000000000001100000000000000111011101001001",
2725 => "0000000000000001000000000000000100000000000000111011101001011",
2726 => "0000000000000001000000000100010100000000000000111011101001101",
2727 => "0000000000000101000000000000001100000000000010011011101001111",
2728 => "0000000000000011000000000000000100000000000000011011101010001",
2729 => "0000000000001011000000000000000100000000000000111011101010100",
2730 => "0000101000001001000000000000000100000000000000011011101010110",
2731 => "0000000000000001000000010010100100000000000000111011101011000",
2732 => "0000000000000101000000000000001100000000000000011011101011010",
2733 => "0000000000000001000000010101000100000000000000111011101011100",
2734 => "0000000000000001000000000000001100000000000000011011101011110",
2735 => "0000000000000001000000000000001100000000000000111011101100000",
2736 => "0000000000000001000000000000001100000000000000011011101100010",
2737 => "0000000000010001000000000000001100000001010000101011101100100",
2738 => "0000000000000001000000000000001100000000010101011011101100110",
2739 => "0000000000000001000000000000001100000000000000111011101101000",
2740 => "0000000000000001000000000000001100000000000000011011101101010",
2741 => "0000000000000001000000000000001100000000000000111011101101100",
2742 => "0000000000000001000000000000000100000000000000111011101101110",
2743 => "0000000000000101000000000000001100000000000000011011101110000",
2744 => "0000000000000001000000000000001100000000000000111011101110010",
2745 => "0000000000101011000000000000001100000000000000011011101110100",
2746 => "0000000000000001000000000000001100000000000000011011101110110",
2747 => "0000000000000011000000000000001100000000000000011011101111000",
2748 => "0000000000000001000000000000001100000000000000011011101111010",
2749 => "0000000000010101000000000000001100000000000000111011101111100",
2750 => "0000000000010101000000000000000100000000000000111011101111110",
2751 => "0000000000000001000000000000001100000000000000111011110000000",
2752 => "0000000000000001000000000000001100000000000000011011110000010",
2753 => "0000000000000001000000100101001000000000000000111011110000100",
2754 => "0000000000000001000000000001000100000000000000011011110000110",
2755 => "0000000000000001000000000000100100000000000000111011110001000",
2756 => "0000000000000001000000000000001100000000100100101011110001010",
2757 => "0000000000000001000000100010000000000000000000111011110001100",
2758 => "0000000000000001000000100101010100000000000000011011110001111",
2759 => "0000000000000001000000000000000100000000000000111011110010001",
2760 => "0000000000000001000000000000001100000000100100101011110010100",
2761 => "0000000000000001000000000000001100000000000000011011110010110",
2762 => "0000000000000001000000000000000100000000000000111011110011000",
2763 => "0000000000000001000000000000001100000000000000111011110011010",
2764 => "0000000000000001000000000000000100000000000000111011110011100",
2765 => "0000000000000001000000000000001100000000000000111011110011110",
2766 => "0000000000000001000000000010000100000000000000111011110100000",
2767 => "0000000000000011000000000000001100000000000000111011110100010",
2768 => "0000000000000101000000000000001100000000010100111011110100100",
2769 => "0000000000000001000000000000001100000000000000111011110100110",
2770 => "0000000000000001000000000100001100000000000000111011110101001",
2771 => "0000000000000011000000000000001100000000001000111011110101100",
2772 => "0000000000000001000000000000001100000000000001011011110101111",
2773 => "0000000100100100000000000000001100000000000000111011110110001",
2774 => "0000000000000001000000101000100000000000000000111011110110011",
2775 => "0000000000000001000000000000001100000000100000101011110110110",
2776 => "0000000000000011000000000000001100000000000000011011110111000",
2777 => "0000000000000001000000000101001100000000000000111011110111011",
2778 => "0000000000000001000000000000000100000000000000011011110111110",
2779 => "0000000000000001000000000001010100000000000000111011111000001",
2780 => "0000000000000011000000000000000100000000000000111011111000100",
2781 => "0000000000000001000000000000001100000000000000111011111000110",
2782 => "0000000000000001000000000000001100000000100000101011111001000",
2783 => "0000000101000001000000000000000100000000000000111011111001010",
2784 => "0000000000000001000000001000000100000000010000001011111001100",
2785 => "0000000100010001000000000000001100000000000001011011111001110",
2786 => "0000000000000001000000000000001100000000000010111011111010000",
2787 => "0000000000101001000000000000001100000000000000111011111010011",
2788 => "0000000000000001000000001010101000000000000000111011111010101",
2789 => "0000010010000101000000000000001100000000000000011011111010111",
2790 => "0000000000000001000000100000101000000000000000101011111011001",
2791 => "0000000000000001000000000000000100000000000000111011111011011",
2792 => "0000001000100010000000000000100100000000000000111011111011101",
2793 => "0000000000000001000000000000001100000000000000011011111011111",
2794 => "0000000000000001000000000000000100000000000000011011111100001",
2795 => "0000000000000001000000000000001100000000100101011011111100100",
2796 => "0000000000000001000000000000001100000000000100011011111100111",
2797 => "0000000000000001000000000000001100000000000000111011111101001",
2798 => "0000000000000001000000000000101100000000000000111011111101100",
2799 => "0000000000000001000000000000100100000000000000111011111101111",
2800 => "0000000000000001000000000001001100000000001010111011111110010",
2801 => "0000000000000001000000000000000100000000000000111011111110101",
2802 => "0000000000000001000000000000001100000000100100101011111111000",
2803 => "0000000000000001000000000001010100000000000000111011111111010",
2804 => "0000000000000011000000000000000100000000000000111011111111100",
2805 => "0000000000000001000000000000001100000000000000111011111111110",
2806 => "0000000000000001000000000000000100000000000000011100000000000",
2807 => "0000000000000001000000000000001100000000000000011100000000010",
2808 => "0000000000000001000000000000001100000000000000011100000000100",
2809 => "0000000001001001000000000000001100000000000000011100000000110",
2810 => "0000000000000001000000000000001100000000000010011100000001000",
2811 => "0000000000000001000000000000000100000000000000111100000001010",
2812 => "0000000010000011000000000000001100000000000000111100000001100",
2813 => "0000000000000001000000000000000100000000000000111100000001110",
2814 => "0000000000001001000000000000001100000000000010011100000010000",
2815 => "0000000000101000000000000000010100000000000000111100000010010",
2816 => "0000000000000001000000000000000100000000000000011100000010100",
2817 => "0000000000000001000000000000001100000000000000111100000010111",
2818 => "0000000000000011000000001001001000000000000000111100000011010",
2819 => "0000000010101011000000000010100100000000000000111100000011100",
2820 => "0000000000000001000000000100010100000000010010011100000011110",
2821 => "0000010000101000000000000000001100000000000000111100000100000",
2822 => "0000000000000001000000000000100100000000000000011100000100010",
2823 => "0000000100010010000000000000001100000000000100011100000100100",
2824 => "0000000000000101000000001010000000000000000000111100000100110",
2825 => "0000000000000001000000000000001100000000000000111100000101000",
2826 => "0000000000000001000000000101010100000000000000011100000101010",
2827 => "0000000010100010000000000000001100000000000100111100000101101",
2828 => "0000000000000001000000010010001000000000000000111100000101111",
2829 => "0000000000000001000000000000001100000000000000111100000110001",
2830 => "0000000000001001000000000000010100000000000000111100000110011",
2831 => "0000000000000001000000000000001100000000000001011100000110101",
2832 => "0000000000000001000000000000000100000000000000111100000110111",
2833 => "0000000000001001000000000000001100000000000000111100000111010",
2834 => "0000000000010011000000000000001100000001000001001100000111100",
2835 => "0000000000000001000000000000000100000000000000111100000111110",
2836 => "0000000000000001000000000000001100000000000010111100001000000",
2837 => "0000000000101000000000000000001100000001001001001100001000010",
2838 => "0000000000000001000000000000001100000000000000011100001000100",
2839 => "0000000000000001000000000000000100000000000000111100001000111",
2840 => "0000000000000001000000000001001100000000000001011100001001001",
2841 => "0000000000000001000000000000001100000000010100011100001001011",
2842 => "0000000000001011000000000000000100000000000000111100001001101",
2843 => "0000000000000011000000000000001100000000000000111100001001111",
2844 => "0000000000000001000000000000000100000000010100101100001010001",
2845 => "0000000000010001000000000000001100000000000000111100001010011",
2846 => "0000000000100011000000001010000000000000000000111100001010101",
2847 => "0000000000100001000000000000001100000000000000111100001011000",
2848 => "0000000000000101000000000000001100000000000000011100001011010",
2849 => "0000000000000001000000000000001100000000000010111100001011100",
2850 => "0000000000000101000000000000001100000001010000101100001011110",
2851 => "0000000001010100000000000000001100000000000000111100001100000",
2852 => "0000000000000011000000000000000100000000000000111100001100011",
2853 => "0000000000000001000000000000010100000000000000111100001100101",
2854 => "0000000000000001000000000000000100000000000010011100001100111",
2855 => "0000000000000001000000000000001100000000000000111100001101001",
2856 => "0000000000000001000000000000001100000000000000011100001101011",
2857 => "0000000000000001000000000000001100000000000100111100001101101",
2858 => "0000000001001011000000000000000000000000001010111100001110000",
2859 => "0000000000100100000000000000001100000000000000111100001110011",
2860 => "0000000000000001000000000000001100000000000000011100001110101",
2861 => "0000000000000001000000000000000100000000000000111100001110111",
2862 => "0000000000000101000000000001000100000000000000111100001111001",
2863 => "0000000000000001000000000001001100000000000000111100001111011",
2864 => "0000010010000011000000000010001000000000000000011100001111101",
2865 => "0000000000000001000000000000001100000000000000011100001111111",
2866 => "0000000000000001000000000000000100000000001010111100010000001",
2867 => "0000000000000001000000000000001100000000000000111100010000100",
2868 => "0000000000000001000000000000001100000000010100011100010000110",
2869 => "0000000000000001000000000000001100000000000000111100010001000",
2870 => "0000000000000001000000000000000100000000000000011100010001010",
2871 => "0000000001001010000000000000001100000000000000111100010001100",
2872 => "0000000100100000000000000010101000000000010101011100010001110",
2873 => "0000000000000001000000000000001100000000000000011100010010000",
2874 => "0000000000100001000000000000000100000000000000111100010010010",
2875 => "0000000000000001000000000000001100000000000000011100010010100",
2876 => "0000000000000001000000000010000100000000000000111100010010111",
2877 => "0000000000001001000000000001000100000000000000111100010011010",
2878 => "0000000000000001000000000000001100000000010010111100010011101",
2879 => "0000000000000011000000000000001100000000000000011100010100000",
2880 => "0000000000000001000000000000101100000000000001011100010100011",
2881 => "0000010100001001000000000000001100000000000000011100010100110",
2882 => "0000000000000001000000000000001100000000000000011100010101001",
2883 => "0000000100100101000000000000001100000000000000111100010101100",
2884 => "0000000000000001000000010010101100000000010100101100010101111",
2885 => "0000000000000001000000000010100100000000000000111100010110001",
2886 => "0000000000000001000000000000001100000000100000001100010110011",
2887 => "0000000010000001000000000000001100000000001000111100010110101",
2888 => "0000000000000001000000001010010100000000000000111100010110111",
2889 => "0000000000000101000000000000001100000000000100111100010111001",
2890 => "0000000000000001000000010000100000000000000000111100010111011",
2891 => "0000000000000001000000000000001100000000000000111100010111101",
2892 => "0000000000000001000000000000001100000000100100101100010111111",
2893 => "0000000000000001000000000000010100000000000000111100011000001",
2894 => "0000000001001010000000000000001100000000000000011100011000011",
2895 => "0000000000000011000000000000001100000001010001011100011000110",
2896 => "0000000000000001000000000000000100000000000000111100011001001",
2897 => "0000000000000001000000000000001100000000000000111100011001011",
2898 => "0000000010000011000000000010001100000000000010111100011001101",
2899 => "0000000000000001000000000000000100000000000000111100011010000",
2900 => "0000000000000001000000000000000100000000000000111100011010011",
2901 => "0000001001001001000000000000001100000000000000111100011010101",
2902 => "0000000000000001000000000000001100000000000000111100011011000",
2903 => "0000000000000001000000000001010100000000000000111100011011010",
2904 => "0000000000000001000000000000001100000000000000111100011011100",
2905 => "0000001000010100000000000000001100000000000000011100011011110",
2906 => "0000000000000001000000000000001100000000000000011100011100000",
2907 => "0000000000000001000000000000001100000000000000111100011100010",
2908 => "0000000000000001000000000000000100000000000000111100011100100",
2909 => "0000000000000001000000000000001100000000000000111100011100110",
2910 => "0000000000000001000000000000001100000000000000011100011101000",
2911 => "0000000000000101000000000000001100000000000000011100011101010",
2912 => "0000000000000001000000000000000100000000000000011100011101100"
);

begin

--process for read and write operation.
PROCESS(clk)
BEGIN
    if(rising_edge(clk)) then
        data_o <= ram(adress);
    end if;
END PROCESS;

end Behavioral;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

--Rectangles--

entity ram_Rectangles is
port ( 	clk : in std_logic;
			adress : in integer;
			data_o : out unsigned(24 downto 0)
     );
end ram_Rectangles;

architecture Behavioral of ram_Rectangles is

--Declaration of type and signal of a 256 element RAM
--with each element being 8 bit wide.
type ram_t is array (0 to 6382) of unsigned(24 downto 0);
signal ram : ram_t := 
(
0 => "0011000100011000100110001",
1 => "0011000111011000001100011",
2 => "0011000100011000011110001",
3 => "0101000100001000011100011",
4 => "0001101001100100100110001",
5 => "0001101100100100001100011",
6 => "0100010010010010011010001",
7 => "0100010100010010001000011",
8 => "0001100101001001001110001",
9 => "0010100101000101001100010",
10 => "0011000101011001000010001",
11 => "0011001101011000100000010",
12 => "0010101000011000011010001",
13 => "0010101011011000001100010",
14 => "0101101110001000101010001",
15 => "0101110011001000010100010",
16 => "0010000000001110011010001",
17 => "0010000011001110001100010",
18 => "0011000110011000011010001",
19 => "0011001000011000001000011",
20 => "0011000100011000011110001",
21 => "0101000100001000011100011",
22 => "0000101000100110110010001",
23 => "0000101100100110010000011",
24 => "0000000010110000001110001",
25 => "0100000010010000001100011",
26 => "0100101001001100111110001",
27 => "0100101110001100010100011",
28 => "0010100110011100101010001",
29 => "0010101011011100010100010",
30 => "0010100000011100100110001",
31 => "0010100011011100001100011",
32 => "0110101011010010011010001",
33 => "1000001011000110011000011",
34 => "0011100101001100101010001",
35 => "0100100101000100101000011",
36 => "0101001000001100101010001",
37 => "0110001000000100101000011",
38 => "0001000101001000100110001",
39 => "0010000101000100100100010",
40 => "1001000000001100101110001",
41 => "1010000000000100101100011",
42 => "0000000110110000110110001",
43 => "0100000110010000110100011",
44 => "0100100110001100100110001",
45 => "0101100110000100100100011",
46 => "0011110010010100011010001",
47 => "0011110100010100001000011",
48 => "0010100111011100110010001",
49 => "0010101101011100011000010",
50 => "0000000011110000001110001",
51 => "0100000011010000001100011",
52 => "0010101000011110011010001",
53 => "0010101011011110001100010",
54 => "0100100110001010111010001",
55 => "0100101101001010011100010",
56 => "0100100101001100101010001",
57 => "0101100101000100101000011",
58 => "0011000110000110110010001",
59 => "0011001100000110011000010",
60 => "0001110101100100001110001",
61 => "0100110101001100001100011",
62 => "0010100110011010011010001",
63 => "0010101000011010001000011",
64 => "1001000001001100111110001",
65 => "1001000001000110111100010",
66 => "0000100001001100111110001",
67 => "0010000001000110111100010",
68 => "0000001000110000111110001",
69 => "0100001000010000111100011",
70 => "0010100110011100110010001",
71 => "0010100110001110011000010",
72 => "0110001100001110011000010",
73 => "0001001100101010110010001",
74 => "0001010000101010010000011",
75 => "0100000001001000101010001",
76 => "0101000001000100101000010",
77 => "0001001101101000101010001",
78 => "0001001101010100101000010",
79 => "0000000001001100110110001",
80 => "0001000001000100110100011",
81 => "1010000010001000110110001",
82 => "1010000010000100110100010",
83 => "0000000101101101001110001",
84 => "0101100101010111001100010",
85 => "1001000100001100100110001",
86 => "1010000100000100100100011",
87 => "0000000011001100101110001",
88 => "0001000011000100101100011",
89 => "0110000001001000100110001",
90 => "0110000001000100100100010",
91 => "0000000110100110001110001",
92 => "0000000111100110000100011",
93 => "0110000001001000100110001",
94 => "0110000001000100100100010",
95 => "0100000001001000100110001",
96 => "0101000001000100100100010",
97 => "0010100101011100111010001",
98 => "0110000101001110011100010",
99 => "0010101100001110011100010",
100 => "0000101010100100001010001",
101 => "0000101011100100000100010",
102 => "1000101101001000101110001",
103 => "1000101101000100101100010",
104 => "0000000100001100100110001",
105 => "0000000111001100001100011",
106 => "0011000100011000100110001",
107 => "0011000111011000001100011",
108 => "0011000101011000011010001",
109 => "0101000101001000011000011",
110 => "0000000001110000010110001",
111 => "0100000001010000010100011",
112 => "0010001010100100011010001",
113 => "0010001100100100001000011",
114 => "0001010001011000011010001",
115 => "0001010001001100001100010",
116 => "0100010100001100001100010",
117 => "1001100011001000110110001",
118 => "1001100011000100110100010",
119 => "0000100011001000110110001",
120 => "0001100011000100110100010",
121 => "0000000001110001011110001",
122 => "0100000001010001011100011",
123 => "0000100111010000110010001",
124 => "0000101011010000010000011",
125 => "0111000111000110111010001",
126 => "0111001110000110011100010",
127 => "0001101100100000011010001",
128 => "0001101100010000001100010",
129 => "0101101111010000001100010",
130 => "0011000110011000011010001",
131 => "0011001000011000001000011",
132 => "0100000111001100110010001",
133 => "0100001101001100011000010",
134 => "0111101111010010011010001",
135 => "0111110001010010001000011",
136 => "0000110001100100001110001",
137 => "0000110010100100000100011",
138 => "0010000100100000110010001",
139 => "0010001010100000011000010",
140 => "0000000001001001010010001",
141 => "0001000001000101010000010",
142 => "0001100000100100001010001",
143 => "0001100001100100000100010",
144 => "0000100101101000111010001",
145 => "0000100101010100011100010",
146 => "0101101100010100011100010",
147 => "0010101000011100110010001",
148 => "0010101100011100010000011",
149 => "0001101110001110100110001",
150 => "0001110001001110001100011",
151 => "0111001111010010011010001",
152 => "0111010001010010001000011",
153 => "0000101111010010011010001",
154 => "0000110001010010001000011",
155 => "0101100110010000101010001",
156 => "0111100110001000010100010",
157 => "0101101011001000010100010",
158 => "0010100101011100111010001",
159 => "0010100101001110011100010",
160 => "0110001100001110011100010",
161 => "0011000000011000010110001",
162 => "0101000000001000010100011",
163 => "0100100000001100100110001",
164 => "0100100011001100001100011",
165 => "0100100110001100100110001",
166 => "0101100110000100100100011",
167 => "0011100000001100100110001",
168 => "0100100000000100100100011",
169 => "0101000110001100100110001",
170 => "0110000110000100100100011",
171 => "0100000110001100100110001",
172 => "0101000110000100100100011",
173 => "0001101000100100010010001",
174 => "0100101000001100010000011",
175 => "0011000000011000100110001",
176 => "0011000011011000001100011",
177 => "0000000000110000011010001",
178 => "0100000000010000011000011",
179 => "0010000111100000110010001",
180 => "0010001011100000010000011",
181 => "0101100110001100011010001",
182 => "0101100110000110011000010",
183 => "0000010100110000001110001",
184 => "0100010100010000001100011",
185 => "0101100110001000100110001",
186 => "0101100110000100100100010",
187 => "0010001101011110010010001",
188 => "0100101101001010010000011",
189 => "0101100110001000100110001",
190 => "0101100110000100100100010",
191 => "0100100110001000100110001",
192 => "0101100110000100100100010",
193 => "0100101100001100110010001",
194 => "0100110010001100011000010",
195 => "0000110110100100001010001",
196 => "0000110111100100000100010",
197 => "0101000111001000101010001",
198 => "0101001100001000010100010",
199 => "0011000111010000101010001",
200 => "0011001100010000010100010",
201 => "0011100110010100011010001",
202 => "0011101000010100001000011",
203 => "0000001110010100010010001",
204 => "0000010000010100001000010",
205 => "0011010010100100001010001",
206 => "0011010011100100000100010",
207 => "0000100001101100001110001",
208 => "0000100010101100000100011",
209 => "0011010000100100001110001",
210 => "0011010001100100000100011",
211 => "0001000100001100111110001",
212 => "0010100100000110111100010",
213 => "1010000100001000101010001",
214 => "1010000100000100101000010",
215 => "0000000100001000101010001",
216 => "0001000100000100101000010",
217 => "0001010000101000011010001",
218 => "0110010000010100001100010",
219 => "0001010011010100001100010",
220 => "0000001100010000100110001",
221 => "0010001100001000100100010",
222 => "0110000000001100100110001",
223 => "0111000000000100100100011",
224 => "0010101010001100011010001",
225 => "0100001010000110011000010",
226 => "0101101000011000011010001",
227 => "1000101000001100001100010",
228 => "0101101011001100001100010",
229 => "0000001000011000011010001",
230 => "0000001000001100001100010",
231 => "0011001011001100001100010",
232 => "0110000000001100100110001",
233 => "0111000000000100100100011",
234 => "0011000000001100100110001",
235 => "0100000000000100100100011",
236 => "0100001110010010011010001",
237 => "0100010000010010001000011",
238 => "0000010000010010011010001",
239 => "0000010010010010001000011",
240 => "0101001000001100101010001",
241 => "0110001000000100101000011",
242 => "0001110011011000001110001",
243 => "0100110011001100001100010",
244 => "0001001010101000001010001",
245 => "0001001011101000000100010",
246 => "0001001001100100110010001",
247 => "0001001001010010011000010",
248 => "0101101111010010011000010",
249 => "0001100000100101100010001",
250 => "0001100000010011100000010",
251 => "0010100110011100101010001",
252 => "0010100110001110010100010",
253 => "0110001011001110010100010",
254 => "0100100101010100110010001",
255 => "0111000101001010011000010",
256 => "0100101011001010011000010",
257 => "0010000101011000110010001",
258 => "0010000101001100011000010",
259 => "0101001011001100011000010",
260 => "0010001110100100001110001",
261 => "0010001111100100000100011",
262 => "0011001101010000100010001",
263 => "0011010001010000010000010",
264 => "0001110000100100011010001",
265 => "0001110011100100001100010",
266 => "0000000000001100011010001",
267 => "0001100000000110011000010",
268 => "0011000110011001001010001",
269 => "0101000110001001001000011",
270 => "0011000001001000111010001",
271 => "0100000001000100111000010",
272 => "0001100010100110001010001",
273 => "0001100011100110000100010",
274 => "0000101000101100110110001",
275 => "0110001000010110110100010",
276 => "0100001001010110010010001",
277 => "0100001011010110001000010",
278 => "0000001100011110101010001",
279 => "0010101100001010101000011",
280 => "0110010000011000011010001",
281 => "1000010000001000011000011",
282 => "0000010000011000011010001",
283 => "0010010000001000011000011",
284 => "1001100001001010110010001",
285 => "1001100101001010010000011",
286 => "0000000010110000010010001",
287 => "0100000010010000010000011",
288 => "0011001000011000010010001",
289 => "0011001010011000001000010",
290 => "0011100101010010011010001",
291 => "0101000101000110011000011",
292 => "0100110001001100011010001",
293 => "0100110100001100001100010",
294 => "0000000111101100111110001",
295 => "0000001100101100010100011",
296 => "0010000001100010100110001",
297 => "0010000100100010001100011",
298 => "0011100101001100101010001",
299 => "0100100101000100101000011",
300 => "1001000001001100100010001",
301 => "1001000001000110100000010",
302 => "0000000001001100011110001",
303 => "0001100001000110011100010",
304 => "1001000000001101011010001",
305 => "1001000000000111011000010",
306 => "0000000000001101011010001",
307 => "0001100000000111011000010",
308 => "1000000111010001000010001",
309 => "1000000111001001000000010",
310 => "0001001010100110011010001",
311 => "0001001100100110001000011",
312 => "0100101001001100110010001",
313 => "0100101101001100010000011",
314 => "0001001111100010011010001",
315 => "0001010001100010001000011",
316 => "0111000111000110111010001",
317 => "0111001110000110011100010",
318 => "0010100110010000101010001",
319 => "0010100110001000010100010",
320 => "0100101011001000010100010",
321 => "0111101000010010101110001",
322 => "1001001000000110101100011",
323 => "0000001000010010101110001",
324 => "0001101000000110101100011",
325 => "0100000110010101001010001",
326 => "0100001111010100100100010",
327 => "0011100111000110111010001",
328 => "0011101110000110011100010",
329 => "0000001110110000100010001",
330 => "0100001110010000100000011",
331 => "0000101010100100111010001",
332 => "0101001010010010111000010",
333 => "0111001100001100011010001",
334 => "0111001111001100001100010",
335 => "0011100000010101000010001",
336 => "0011100000001010100000010",
337 => "0110001000001010100000010",
338 => "0101000000010010011010001",
339 => "0110100000000110011000011",
340 => "0010000011100000010010001",
341 => "0110000011010000010000010",
342 => "0101000000010010011010001",
343 => "0110100000000110011000011",
344 => "0000100001101000010010001",
345 => "0000100001010100001000010",
346 => "0101100011010100001000010",
347 => "0101000000010010011010001",
348 => "0110100000000110011000011",
349 => "0010100000010010011010001",
350 => "0100000000000110011000011",
351 => "0100010010010100011010001",
352 => "0100010100010100001000011",
353 => "0011000011001100100110001",
354 => "0100000011000100100100011",
355 => "0011100011011000011010001",
356 => "0011100101011000001000011",
357 => "0000001010100100001110001",
358 => "0000001011100100000100011",
359 => "0000101010101100001110001",
360 => "0000101011101100000100011",
361 => "0010101011010000100010001",
362 => "0100101011001000100000010",
363 => "0110001011001100011010001",
364 => "0110001011000110011000010",
365 => "0011001011001100011010001",
366 => "0100101011000110011000010",
367 => "0011101010010110011010001",
368 => "0011101100010110001000011",
369 => "0000001101110000010010001",
370 => "0000001101011000001000010",
371 => "0110001111011000001000010",
372 => "0001000100101100110010001",
373 => "0110100100010110011000010",
374 => "0001001010010110011000010",
375 => "0001000000101001000110001",
376 => "0110000000010101000100010",
377 => "0111000000000101100010001",
378 => "0111000000000011100000010",
379 => "0100000000000101100010001",
380 => "0100100000000011100000010",
381 => "0111000001000101011010001",
382 => "0111000001000011011000010",
383 => "0100000001000101011010001",
384 => "0100100001000011011000010",
385 => "1000100110000111001010001",
386 => "1001000110000011001000011",
387 => "0011001110010010011010001",
388 => "0011010000010010001000011",
389 => "0110101110010010010010001",
390 => "0110110000010010001000010",
391 => "0001110010100100001110001",
392 => "0001110011100100000100011",
393 => "0100100100010001001010001",
394 => "0110100100001000100100010",
395 => "0100101101001000100100010",
396 => "0000010001100100001110001",
397 => "0000010010100100000100011",
398 => "0000000010011000010010001",
399 => "0011000010001100010000010",
400 => "0011001000011100011010001",
401 => "0011001011011100001100010",
402 => "0011100101001100011010001",
403 => "0101000101000110011000010",
404 => "0101000101001101000010001",
405 => "0101001101001100100000010",
406 => "0000100100010011000010001",
407 => "0010000100000111000000011",
408 => "0010100000100100100110001",
409 => "0010100011100100001100011",
410 => "0100101111001010100010001",
411 => "0100110011001010010000010",
412 => "1010000000001000100110001",
413 => "1010000000000100100100010",
414 => "0001000000100100001110001",
415 => "0001000001100100000100011",
416 => "0010110110100110001010001",
417 => "0010110111100110000100010",
418 => "0000000000001000100110001",
419 => "0001000000000100100100010",
420 => "0010100110100111001010001",
421 => "0010101100100110011000011",
422 => "0000000001001100100110001",
423 => "0001000001000100100100011",
424 => "0011000101011100110010001",
425 => "0110100101001110011000010",
426 => "0011001011001110011000010",
427 => "0000000001101000001010001",
428 => "0000000010101000000100010",
429 => "0000100010101100001110001",
430 => "0000100011101100000100011",
431 => "0001001000001110100110001",
432 => "0001001011001110001100011",
433 => "0001001100101100010010001",
434 => "0110101100010110001000010",
435 => "0001001110010110001000010",
436 => "0000001100101100010010001",
437 => "0000001100010110001000010",
438 => "0101101110010110001000010",
439 => "0100100111001100101110001",
440 => "0101100111000100101100011",
441 => "0011100001010010011010001",
442 => "0101000001000110011000011",
443 => "0101100010001000101010001",
444 => "0101100111001000010100010",
445 => "0011000100011000110010001",
446 => "0011001010011000011000010",
447 => "1001000001001100111110001",
448 => "1001000110001100010100011",
449 => "0001101111100100001110001",
450 => "0001110000100100000100011",
451 => "1001000101001100100110001",
452 => "1001001000001100001100011",
453 => "0000100101100000011010001",
454 => "0000100101010000001100010",
455 => "0100101000010000001100010",
456 => "0101100000001100100110001",
457 => "0110100000000100100100011",
458 => "0000000100110000111010001",
459 => "0000000100011000011100010",
460 => "0110001011011000011100010",
461 => "0110100000001000110110001",
462 => "0110100000000100110100010",
463 => "0011100000001000110110001",
464 => "0100100000000100110100010",
465 => "0101100110001100100110001",
466 => "0110100110000100100100011",
467 => "0100000111001100100110001",
468 => "0101000111000100100100011",
469 => "0110110001010010011010001",
470 => "0110110011010010001000011",
471 => "0001010010011100011010001",
472 => "0001010010001110001100010",
473 => "0100110101001110001100010",
474 => "0001110010100100010010001",
475 => "0110010010010010001000010",
476 => "0001110100010010001000010",
477 => "0000010100011110010010001",
478 => "0010110100001010010000011",
479 => "0100101111011110100110001",
480 => "0111001111001010100100011",
481 => "0010000100100000010010001",
482 => "0010000110100000001000010",
483 => "0011100110010100011010001",
484 => "0011101000010100001000011",
485 => "0000001110011110101010001",
486 => "0010101110001010101000011",
487 => "0011101001010100111010001",
488 => "0110001001001010011100010",
489 => "0011110000001010011100010",
490 => "0011100110001100100110001",
491 => "0100100110000100100100011",
492 => "0001100110100100001110001",
493 => "0001100111100100000100011",
494 => "0000001010100100001110001",
495 => "0000001011100100000100011",
496 => "0001110000100100010010001",
497 => "0110010000010010001000010",
498 => "0001110010010010001000010",
499 => "0010000110011100011010001",
500 => "0010000110001110001100010",
501 => "0101101001001110001100010",
502 => "0110100000000101001010001",
503 => "0110100000000011001000010",
504 => "0100100000000101001010001",
505 => "0101000000000011001000010",
506 => "0010100111011110101010001",
507 => "0101000111001010101000011",
508 => "0000110100101010010010001",
509 => "0100010100001110010000011",
510 => "0101000101001011001010001",
511 => "0101001110001010100100010",
512 => "0000000010110000011010001",
513 => "0000000010011000001100010",
514 => "0110000101011000001100010",
515 => "0000100001101100100010001",
516 => "0110000001010110010000010",
517 => "0000100101010110010000010",
518 => "0010000000011110100110001",
519 => "0010000011011110001100011",
520 => "0000000000110001001110001",
521 => "0100000000010001001100011",
522 => "0001010101100100001110001",
523 => "0101110101010010001100010",
524 => "0100100111010100010010001",
525 => "0100100111001010010000010",
526 => "0010100111010100010010001",
527 => "0101000111001010010000010",
528 => "1000101000001101000010001",
529 => "1010001000000110100000010",
530 => "1000110000000110100000010",
531 => "0000101111101000010010001",
532 => "0000101111010100001000010",
533 => "0101110001010100001000010",
534 => "0111001111010100011010001",
535 => "0111010001010100001000011",
536 => "0001100000100000100110001",
537 => "0001100011100000001100011",
538 => "0111100110001110111110001",
539 => "0111101011001110010100011",
540 => "0100100001001100110110001",
541 => "0101100001000100110100011",
542 => "1000100010001100111010001",
543 => "1000100010000110111000010",
544 => "0001101110011000101010001",
545 => "0001101110001100010100010",
546 => "0100110011001100010100010",
547 => "0011100110010100011010001",
548 => "0011101000010100001000011",
549 => "0000100010001100111010001",
550 => "0010000010000110111000010",
551 => "0101000100001010110010001",
552 => "0101001000001010010000011",
553 => "0000010001110000010110001",
554 => "0100010001010000010100011",
555 => "0111100111001010110010001",
556 => "0111101011001010010000011",
557 => "0001100001001100110010001",
558 => "0001100001000110011000010",
559 => "0011000111000110011000010",
560 => "0110001101001100011010001",
561 => "0110010000001100001100010",
562 => "0011001101001100011010001",
563 => "0011010000001100001100010",
564 => "0111000110000111000010001",
565 => "0111001110000110100000010",
566 => "0000101100011010011010001",
567 => "0000101110011010001000011",
568 => "0110100001001000100110001",
569 => "0110100001000100100100010",
570 => "0011100000010010011010001",
571 => "0101000000000110011000011",
572 => "0110000010001100100110001",
573 => "0110000010000110100100010",
574 => "0011000010001100100110001",
575 => "0100100010000110100100010",
576 => "0011010010011000011010001",
577 => "0011010100011000001000011",
578 => "0011100110001100100110001",
579 => "0100100110000100100100011",
580 => "0011100111011000001110001",
581 => "0011100111001100001100010",
582 => "0100000011010001010110001",
583 => "0100001010010000011100011",
584 => "0011100100010100110010001",
585 => "0011101000010100010000011",
586 => "0000000001001100100110001",
587 => "0000000100001100001100011",
588 => "0111100010000101010010001",
589 => "0111100010000011010000010",
590 => "0000000011001100100110001",
591 => "0000000110001100001100011",
592 => "0111100011000101010110001",
593 => "0111100011000011010100010",
594 => "0011100000000101011110001",
595 => "0100000000000011011100010",
596 => "0111101000010010010010001",
597 => "0111101010010010001000010",
598 => "0000001000010010010010001",
599 => "0000001010010010001000010",
600 => "0100001110010010011010001",
601 => "0100010000010010001000011",
602 => "0000001110010010011010001",
603 => "0000010000010010001000011",
604 => "0001101010100100010010001",
605 => "0100101010001100010000011",
606 => "0000000000110001001110001",
607 => "0100000000010001001100011",
608 => "0100100001010000110010001",
609 => "0100100111010000011000010",
610 => "0101000110001000101010001",
611 => "0110000110000100101000010",
612 => "0011101001010100110010001",
613 => "0110001001001010011000010",
614 => "0011101111001010011000010",
615 => "0010100000000111001110001",
616 => "0011000000000011001100011",
617 => "0111000000001100101010001",
618 => "1000000000000100101000011",
619 => "0001000000001100110010001",
620 => "0001000000000110011000010",
621 => "0010100110000110011000010",
622 => "0000001011110000001010001",
623 => "0000001100110000000100010",
624 => "0010001001011010010010001",
625 => "0010001011011010001000010",
626 => "0100101000001100100110001",
627 => "0100101011001100001100011",
628 => "0000001100100000010010001",
629 => "0000001110100000001000010",
630 => "1001001100001100100110001",
631 => "1001001111001100001100011",
632 => "0000001100001100100110001",
633 => "0000001111001100001100011",
634 => "0100000111010100010010001",
635 => "0100000111001010010000010",
636 => "0100000111001100100110001",
637 => "0101000111000100100100011",
638 => "0101100000001100100110001",
639 => "0110100000000100100100011",
640 => "0011100000001100100110001",
641 => "0100100000000100100100011",
642 => "0110000011001100111110001",
643 => "0111000011000100111100011",
644 => "0011000011001100111110001",
645 => "0100000011000100111100011",
646 => "0111100010010010010010001",
647 => "0111100100010010001000010",
648 => "0010101010001100011110001",
649 => "0100001010000110011100010",
650 => "0100101110001100101010001",
651 => "0100110011001100010100010",
652 => "0011101101001010100010001",
653 => "0011110001001010010000010",
654 => "0111000101000111000010001",
655 => "0111001101000110100000010",
656 => "0001010001100100001110001",
657 => "0001010010100100000100011",
658 => "0010110010100110001110001",
659 => "0010110011100110000100011",
660 => "0100100000001100100110001",
661 => "0101100000000100100100011",
662 => "0110000100000111001010001",
663 => "0110100100000011001000011",
664 => "0100100100000111001010001",
665 => "0101000100000011001000011",
666 => "0001100011100100100110001",
667 => "0100100011001100100100011",
668 => "0011000001001100111010001",
669 => "0100000001000100111000011",
670 => "0110010000010010011010001",
671 => "0110010011010010001100010",
672 => "0000100011101001000010001",
673 => "0000100011010100100000010",
674 => "0101101011010100100000010",
675 => "0110000101001100110010001",
676 => "0111100101000110011000010",
677 => "0110001011000110011000010",
678 => "0000100010101101000010001",
679 => "0000100010010110100000010",
680 => "0110001010010110100000010",
681 => "0101001110001010101010001",
682 => "0101010011001010010100010",
683 => "0001110101100100001110001",
684 => "0001110110100100000100011",
685 => "0101001110001100101010001",
686 => "0110001110000100101000011",
687 => "0000000010110000010010001",
688 => "0100000010010000010000011",
689 => "0011000100011000100110001",
690 => "0011000111011000001100011",
691 => "0011000110011000010110001",
692 => "0101000110001000010100011",
693 => "0010101000011100110010001",
694 => "0010101100011100010000011",
695 => "0010001110010000101010001",
696 => "0010001110001000010100010",
697 => "0100010011001000010100010",
698 => "0101100110001010111010001",
699 => "0101101101001010011100010",
700 => "0011100110000111000010001",
701 => "0011101110000110100000010",
702 => "0001100111100100100010001",
703 => "0100100111001100100000011",
704 => "0001000011101000001010001",
705 => "0001000100101000000100010",
706 => "0001101100100110011010001",
707 => "0001101110100110001000011",
708 => "0100000110001100100110001",
709 => "0101000110000100100100011",
710 => "1000000110001100111010001",
711 => "1000000110000110111000010",
712 => "0011101001001100110010001",
713 => "0100101001000100110000011",
714 => "1001000110001101001010001",
715 => "1010100110000110100100010",
716 => "1001001111000110100100010",
717 => "0000000110001101001010001",
718 => "0000000110000110100100010",
719 => "0001101111000110100100010",
720 => "1001000010001100100110001",
721 => "1001000101001100001100011",
722 => "0001110010011110011010001",
723 => "0001110100011110001000011",
724 => "1001000010001100100110001",
725 => "1001000101001100001100011",
726 => "0000000010001100100110001",
727 => "0000000101001100001100011",
728 => "0010101010100100001010001",
729 => "0010101011100100000100010",
730 => "0011000000011000011010001",
731 => "0011000010011000001000011",
732 => "0101000000001100100110001",
733 => "0110000000000100100100011",
734 => "0100000000001100100110001",
735 => "0101000000000100100100011",
736 => "0111101100010010011010001",
737 => "0111101110010010001000011",
738 => "0001100110011010011010001",
739 => "0001101000011010001000011",
740 => "0111101100010010011010001",
741 => "0111101110010010001000011",
742 => "0001000101001100111110001",
743 => "0010100101000110111100010",
744 => "0100001000010010011010001",
745 => "0101101000000110011000011",
746 => "0100000110000110111010001",
747 => "0100001101000110011100010",
748 => "0111101100010010011010001",
749 => "0111101110010010001000011",
750 => "0010001100010100010010001",
751 => "0100101100001010010000010",
752 => "0110100001001001001110001",
753 => "0110100001000101001100010",
754 => "0011100001001001001110001",
755 => "0100100001000101001100010",
756 => "1001001001001100100110001",
757 => "1001001100001100001100011",
758 => "0000110101100100001110001",
759 => "0000110110100100000100011",
760 => "0111001101010100100110001",
761 => "0111010000010100001100011",
762 => "0000101101101100010010001",
763 => "0000101101010110001000010",
764 => "0110001111010110001000010",
765 => "0010000110100000011010001",
766 => "0110000110010000001100010",
767 => "0010001001010000001100010",
768 => "0000100000100101011010001",
769 => "0000100000010010101100010",
770 => "0101001011010010101100010",
771 => "0101000111010000111010001",
772 => "0111000111001000011100010",
773 => "0101001110001000011100010",
774 => "0000000100001101010010001",
775 => "0000000100000110101000010",
776 => "0001101110000110101000010",
777 => "0111100000001100100110001",
778 => "1000100000000100100100011",
779 => "0001100000001100100110001",
780 => "0010100000000100100100011",
781 => "0111101100001100110010001",
782 => "1001001100000110011000010",
783 => "0111110010000110011000010",
784 => "0001101100001100110010001",
785 => "0001101100000110011000010",
786 => "0011010010000110011000010",
787 => "0111101100010010011010001",
788 => "0111101110010010001000011",
789 => "0000001100010010011010001",
790 => "0000001110010010001000011",
791 => "0010001110100110001110001",
792 => "0010001111100110000100011",
793 => "0001001101100110001110001",
794 => "0001001110100110000100011",
795 => "0111001111010100011010001",
796 => "0111010001010100001000011",
797 => "0011000000010100110010001",
798 => "0011000000001010011000010",
799 => "0101100110001010011000010",
800 => "1000100001001100110010001",
801 => "1010000001000110011000010",
802 => "1000100111000110011000010",
803 => "0000100001001100110010001",
804 => "0000100001000110011000010",
805 => "0010000111000110011000010",
806 => "1000001110001100100110001",
807 => "1000010001001100001100011",
808 => "0011100011010010110010001",
809 => "0011101001010010011000010",
810 => "0110000001001000110010001",
811 => "0110000111001000011000010",
812 => "0010000000011100100010001",
813 => "0010000100011100010000010",
814 => "0101000110001100100110001",
815 => "0110000110000100100100011",
816 => "0001001010100100001110001",
817 => "0100001010001100001100011",
818 => "0111101111010010011010001",
819 => "0111110001010010001000011",
820 => "0000000001101011011110001",
821 => "0011100001001111011100011",
822 => "0011001001100010010010001",
823 => "0011001011100010001000010",
824 => "0000100000010111001010001",
825 => "0000100110010110011000011",
826 => "0011001111011010011010001",
827 => "0011010001011010001000011",
828 => "0000001111010010011010001",
829 => "0000010001010010001000011",
830 => "0100000111011110010010001",
831 => "0110100111001010010000011",
832 => "0100101100001100100110001",
833 => "0100101111001100001100011",
834 => "0011001000100100001110001",
835 => "0110001000001100001100011",
836 => "0000001110110000010010001",
837 => "0100001110010000010000011",
838 => "1000001010000110110010001",
839 => "1000010000000110011000010",
840 => "0000000011110000001110001",
841 => "0000000100110000000100011",
842 => "0111010001010100011010001",
843 => "0111010011010100001000011",
844 => "0000101101100100001110001",
845 => "0011101101001100001100011",
846 => "0010100000100100100110001",
847 => "0010100011100100001100011",
848 => "0010000011100000100110001",
849 => "0010000110100000001100011",
850 => "1000000101000110110010001",
851 => "1000001011000110011000010",
852 => "0000000111100100010010001",
853 => "0011000111001100010000011",
854 => "0101000110001100100110001",
855 => "0110000110000100100100011",
856 => "0100101000001100101010001",
857 => "0101101000000100101000011",
858 => "0100101111001100100110001",
859 => "0101101111000100100100011",
860 => "0001100001100101010110001",
861 => "0110000001010011010100010",
862 => "0011001000011000011110001",
863 => "0011001000001100011100010",
864 => "0100000101001100100110001",
865 => "0101000101000100100100011",
866 => "0000000010110000010010001",
867 => "0100000010010000010000011",
868 => "0111000111001010110010001",
869 => "0111001011001010010000011",
870 => "0010100111001010110010001",
871 => "0010101011001010010000011",
872 => "0100100110001100100110001",
873 => "0101100110000100100100011",
874 => "0000000001001101000110001",
875 => "0001100001000111000100010",
876 => "0001100001100110100110001",
877 => "0001100100100110001100011",
878 => "0001110010011000011010001",
879 => "0001110010001100001100010",
880 => "0100110101001100001100010",
881 => "1010000100001001001110001",
882 => "1010000100000101001100010",
883 => "0000010000010100011110001",
884 => "0010110000001010011100010",
885 => "0100000111010100110010001",
886 => "0110100111001010011000010",
887 => "0100001101001010011000010",
888 => "0011000111010100110010001",
889 => "0011000111001010011000010",
890 => "0101101101001010011000010",
891 => "0100100010010010011010001",
892 => "0110000010000110011000011",
893 => "0000110100101010010010001",
894 => "0100010100001110010000011",
895 => "0100101100010010011010001",
896 => "0100101110010010001000011",
897 => "0011100010010010011010001",
898 => "0101000010000110011000011",
899 => "0110100000001000111010001",
900 => "0110100000000100111000010",
901 => "0011100000001000111010001",
902 => "0100100000000100111000010",
903 => "0111001111010010011010001",
904 => "0111010001010010001000011",
905 => "0001001000100100010110001",
906 => "0100001000001100010100011",
907 => "1001000011001100101110001",
908 => "1010000011000100101100011",
909 => "0011000101010110111010001",
910 => "0011001100010110011100010",
911 => "1001000100001100100110001",
912 => "1001000111001100001100011",
913 => "0011100110010010011010001",
914 => "0011101000010010001000011",
915 => "1001000100001100100110001",
916 => "1001000111001100001100011",
917 => "0000000100001100100110001",
918 => "0000000111001100001100011",
919 => "0100100100010010010010001",
920 => "0100100110010010001000010",
921 => "0000010110100110001010001",
922 => "0000010111100110000100010",
923 => "1000101110001100100110001",
924 => "1000110001001100001100011",
925 => "0000101110001100100110001",
926 => "0000110001001100001100011",
927 => "0111001011001000100110001",
928 => "0111001011000100100100010",
929 => "0011001011001000100110001",
930 => "0100001011000100100100010",
931 => "0001101001100100011110001",
932 => "0100101001001100011100011",
933 => "0100101100001100101010001",
934 => "0100110001001100010100010",
935 => "0110000000001100100110001",
936 => "0111000000000100100100011",
937 => "0011000000001100100110001",
938 => "0100000000000100100100011",
939 => "0011010001100100001110001",
940 => "0011010010100100000100011",
941 => "0000110001100100001110001",
942 => "0000110010100100000100011",
943 => "0101000110010110110010001",
944 => "0101001100010110011000010",
945 => "0010100110011100011010001",
946 => "0010100110001110001100010",
947 => "0110001001001110001100010",
948 => "0010100100011110010010001",
949 => "0010100110011110001000010",
950 => "0000000000101100001010001",
951 => "0000000001101100000100010",
952 => "0000000000110001100010001",
953 => "0100000000010001100000011",
954 => "0000101111100100010010001",
955 => "0101001111010010010000010",
956 => "0011001000011000100110001",
957 => "0011001011011000001100011",
958 => "0010001100001110110010001",
959 => "0010010000001110010000011",
960 => "0000100010101100011010001",
961 => "0110000010010110001100010",
962 => "0000100101010110001100010",
963 => "0010110100011100001110001",
964 => "0110010100001110001100010",
965 => "0000000000110001000010001",
966 => "0110000000011000100000010",
967 => "0000001000011000100000010",
968 => "0001101101100100010010001",
969 => "0001101101010010001000010",
970 => "0110001111010010001000010",
971 => "0001001010101100001010001",
972 => "0001001011101100000100010",
973 => "0011000011010110100010001",
974 => "0011000111010110010000010",
975 => "0111000101001100011010001",
976 => "0111001000001100001100010",
977 => "0000000111110000011010001",
978 => "0000001001110000001000011",
979 => "0111000000010100101010001",
980 => "1001100000001010010100010",
981 => "0111000101001010010100010",
982 => "0000000000010100101010001",
983 => "0000000000001010010100010",
984 => "0010100101001010010100010",
985 => "0000000001110000010010001",
986 => "0110000001011000001000010",
987 => "0000000011011000001000010",
988 => "0000010001100100001110001",
989 => "0000010010100100000100011",
990 => "0010101111100000011010001",
991 => "0110101111010000001100010",
992 => "0010110010010000001100010",
993 => "0001101111100000011010001",
994 => "0001101111010000001100010",
995 => "0101110010010000001100010",
996 => "0011010000100100001110001",
997 => "0011010001100100000100011",
998 => "0000001101101010101010001",
999 => "0000010010101010010100010",
1000 => "0110100000001101100010001",
1001 => "0111100000000101100000011",
1002 => "0011100100001100101110001",
1003 => "0100100100000100101100011",
1004 => "0100100101010010011010001",
1005 => "0110000101000110011000011",
1006 => "0000100100000101010010001",
1007 => "0000101110000100101000010",
1008 => "0110100000001101100010001",
1009 => "0111100000000101100000011",
1010 => "0010100000001101100010001",
1011 => "0011100000000101100000011",
1012 => "1000000111001100111010001",
1013 => "1001100111000110011100010",
1014 => "1000001110000110011100010",
1015 => "0010000111001000110010001",
1016 => "0011000111000100110000010",
1017 => "0000000101110000111010001",
1018 => "0100000101010000111000011",
1019 => "0010101101010100011010001",
1020 => "0010101111010100001000011",
1021 => "0110000000001100100110001",
1022 => "0111000000000100100100011",
1023 => "0001000111001100111010001",
1024 => "0001000111000110011100010",
1025 => "0010101110000110011100010",
1026 => "0111100010010010111110001",
1027 => "1001000010000110111100011",
1028 => "0000000010001100100110001",
1029 => "0001000010000100100100011",
1030 => "0110000010010100111010001",
1031 => "1000100010001010011100010",
1032 => "0110001001001010011100010",
1033 => "0101100110000101001010001",
1034 => "0110000110000011001000010",
1035 => "0100100101011110011010001",
1036 => "0111000101001010011000011",
1037 => "0100000110001100101010001",
1038 => "0101000110000100101000011",
1039 => "0110000000001100100110001",
1040 => "0111000000000100100100011",
1041 => "0001100011010010011110001",
1042 => "0011000011000110011100011",
1043 => "0011000111011100001110001",
1044 => "0011000111001110001100010",
1045 => "0011100111010000011010001",
1046 => "0101100111001000011000010",
1047 => "0110000111001110110010001",
1048 => "0110001101001110011000010",
1049 => "0101000110001001001010001",
1050 => "0101000110000100100100010",
1051 => "0110001111000100100100010",
1052 => "1000001110001100100110001",
1053 => "1000010001001100001100011",
1054 => "0010000000001100110110001",
1055 => "0011000000000100110100011",
1056 => "0001000010101010001110001",
1057 => "0100100010001110001100011",
1058 => "0010100100001010110010001",
1059 => "0010101000001010010000011",
1060 => "0101000011001000101010001",
1061 => "0101001000001000010100010",
1062 => "0100000100001010100010001",
1063 => "0100001000001010010000010",
1064 => "0011000000010110100110001",
1065 => "0011000011010110001100011",
1066 => "0011000110011000010110001",
1067 => "0101000110001000010100011",
1068 => "0000000000110000010110001",
1069 => "0100000000010000010100011",
1070 => "0000101010101110011010001",
1071 => "0000101100101110001000011",
1072 => "0001110101100100001110001",
1073 => "0100110101001100001100011",
1074 => "0001100110101010011010001",
1075 => "0001101000101010001000011",
1076 => "0000000101001100110010001",
1077 => "0001000101000100110000011",
1078 => "0101000010001000111110001",
1079 => "0101000111001000010100011",
1080 => "0100000111010000101010001",
1081 => "0100001100010000010100010",
1082 => "0010100111011110110010001",
1083 => "0101000111001010110000011",
1084 => "0000010001010100011010001",
1085 => "0000010011010100001000011",
1086 => "0111010010010010011010001",
1087 => "0111010100010010001000011",
1088 => "0100100110001101000010001",
1089 => "0100101110001100100000010",
1090 => "0111010010010010011010001",
1091 => "0111010100010010001000011",
1092 => "0000110010010010011010001",
1093 => "0000110100010010001000011",
1094 => "0111101001010010011010001",
1095 => "0111101011010010001000011",
1096 => "0000001001010010011010001",
1097 => "0000001011010010001000011",
1098 => "1000100011001100100110001",
1099 => "1001100011000100100100011",
1100 => "0001010001100100001110001",
1101 => "0001010010100100000100011",
1102 => "0001101111101010011010001",
1103 => "0001110001101010001000011",
1104 => "0100110001001100011010001",
1105 => "0100110100001100001100010",
1106 => "1001000011001100100110001",
1107 => "1001000110001100001100011",
1108 => "0000000011001100100110001",
1109 => "0000000110001100001100011",
1110 => "0010000000100000101010001",
1111 => "0110000000010000010100010",
1112 => "0010000101010000010100010",
1113 => "0001000000010101000010001",
1114 => "0001000000001010100000010",
1115 => "0011101000001010100000010",
1116 => "0111000000010100010110001",
1117 => "0111000000001010010100010",
1118 => "0000000000010100010110001",
1119 => "0010100000001010010100010",
1120 => "1001000011001100101010001",
1121 => "1001000011000110101000010",
1122 => "0010101011011000011010001",
1123 => "0010101011001100001100010",
1124 => "0101101110001100001100010",
1125 => "1010100000000111001010001",
1126 => "1011000000000011001000011",
1127 => "0011000000001100100110001",
1128 => "0100000000000100100100011",
1129 => "0100001000010010011110001",
1130 => "0101101000000110011100011",
1131 => "0011101100010000101010001",
1132 => "0011101100001000010100010",
1133 => "0101110001001000010100010",
1134 => "1010100000000111001010001",
1135 => "1011000000000011001000011",
1136 => "0101000110001000100110001",
1137 => "0110000110000100100100010",
1138 => "0111100000010010011010001",
1139 => "0111100010010010001000011",
1140 => "0000000010110000001110001",
1141 => "0000000011110000000100011",
1142 => "0101100111001100100110001",
1143 => "0110100111000100100100011",
1144 => "0011100110001100101010001",
1145 => "0100100110000100101000011",
1146 => "0110000001001100110010001",
1147 => "0111000001000100110000011",
1148 => "0011000100011000110010001",
1149 => "0011001010011000011000010",
1150 => "0111000011000101010110001",
1151 => "0111000011000011010100010",
1152 => "0011000001011000100010001",
1153 => "0011000101011000010000010",
1154 => "0001100000100100100010001",
1155 => "0001100100100100010000010",
1156 => "0001100000100100001110001",
1157 => "0001100001100100000100011",
1158 => "0000001101110000010010001",
1159 => "0110001101011000001000010",
1160 => "0000001111011000001000010",
1161 => "0101000101001000100110001",
1162 => "0110000101000100100100010",
1163 => "0101100001001100100110001",
1164 => "0110100001000100100100011",
1165 => "0011000010001101011010001",
1166 => "0100000010000101011000011",
1167 => "1000001010010000111010001",
1168 => "1010001010001000011100010",
1169 => "1000010001001000011100010",
1170 => "0001100100100000111110001",
1171 => "0001101001100000010100011",
1172 => "1000001010010000111010001",
1173 => "1010001010001000011100010",
1174 => "1000010001001000011100010",
1175 => "0000001010010000111010001",
1176 => "0000001010001000011100010",
1177 => "0010010001001000011100010",
1178 => "0101001110010110011010001",
1179 => "0101010001010110001100010",
1180 => "0000000111110000100110001",
1181 => "0100000111010000100100011",
1182 => "0110100001001001000010001",
1183 => "0110100001000101000000010",
1184 => "0011100001001001000010001",
1185 => "0100100001000101000000010",
1186 => "0010100101100000100010001",
1187 => "0110100101010000010000010",
1188 => "0010101001010000010000010",
1189 => "0000001001001100100110001",
1190 => "0000001100001100001100011",
1191 => "0011010000100100001110001",
1192 => "0011010001100100000100011",
1193 => "0001101100001100100110001",
1194 => "0001101111001100001100011",
1195 => "0100001110010010011010001",
1196 => "0100010000010010001000011",
1197 => "0001001101010000101010001",
1198 => "0001001101001000010100010",
1199 => "0011010010001000010100010",
1200 => "0111100101000111001010001",
1201 => "0111101011000110011000011",
1202 => "0001100101100100001110001",
1203 => "0001100110100100000100011",
1204 => "1000100101001100101110001",
1205 => "1001100101000100101100011",
1206 => "0000100101001100101110001",
1207 => "0001100101000100101100011",
1208 => "1001100001001000100110001",
1209 => "1001100001000100100100010",
1210 => "0000100001001000100110001",
1211 => "0001100001000100100100010",
1212 => "0010001111100100100110001",
1213 => "0010001111010010100100010",
1214 => "0011001001011000010010001",
1215 => "0011001011011000001000010",
1216 => "0111100010010010011010001",
1217 => "0111100100010010001000011",
1218 => "0000000010010010011010001",
1219 => "0000000100010010001000011",
1220 => "0111100000001101000110001",
1221 => "1000100000000101000100011",
1222 => "0001100000001101000110001",
1223 => "0010100000000101000100011",
1224 => "0100010001010010010010001",
1225 => "0100010011010010001000010",
1226 => "0011000101000111001010001",
1227 => "0011001011000110011000011",
1228 => "0010100010011100110010001",
1229 => "0010101000011100011000010",
1230 => "0101000010000110110010001",
1231 => "0101001000000110011000010",
1232 => "0101000111011100111110001",
1233 => "0101001100011100010100011",
1234 => "0000000111011100111110001",
1235 => "0000001100011100010100011",
1236 => "0111100000010010011010001",
1237 => "0111100010010010001000011",
1238 => "0000000000010010011010001",
1239 => "0000000010010010001000011",
1240 => "0110000110001100111010001",
1241 => "0111000110000100111000011",
1242 => "0100100111001100100110001",
1243 => "0101100111000100100100011",
1244 => "0110000110001100111110001",
1245 => "0111000110000100111100011",
1246 => "0011000110001100111110001",
1247 => "0100000110000100111100011",
1248 => "0111100011010000100110001",
1249 => "0111100011001000100100010",
1250 => "0000000000010011010110001",
1251 => "0001100000000111010100011",
1252 => "0101101001010000110010001",
1253 => "0101101101010000010000011",
1254 => "0011000111010100110010001",
1255 => "0011000111001010011000010",
1256 => "0101101101001010011000010",
1257 => "0101000110001001001010001",
1258 => "0110000110000100100100010",
1259 => "0101001111000100100100010",
1260 => "0000000000001100100110001",
1261 => "0000000011001100001100011",
1262 => "0001101110100100001110001",
1263 => "0001101111100100000100011",
1264 => "0001101110010000101010001",
1265 => "0001101110001000010100010",
1266 => "0011110011001000010100010",
1267 => "0000001100110000010010001",
1268 => "0110001100011000001000010",
1269 => "0000001110011000001000010",
1270 => "0000000010000111010010001",
1271 => "0000100010000011010000011",
1272 => "0110010000010100100010001",
1273 => "1000110000001010010000010",
1274 => "0110010100001010010000010",
1275 => "0001010000010100100010001",
1276 => "0001010000001010010000010",
1277 => "0011110100001010010000010",
1278 => "0011100000010100100110001",
1279 => "0011100011010100001100011",
1280 => "0000000000110000001110001",
1281 => "0100000000010000001100011",
1282 => "0001101000011110010010001",
1283 => "0001101010011110001000010",
1284 => "0011000101011000011010001",
1285 => "0101000101001000011000011",
1286 => "0010101101011100011010001",
1287 => "0010110000011100001100010",
1288 => "0101101110001000101010001",
1289 => "0101110011001000010100010",
1290 => "0000000110001100011110001",
1291 => "0001100110000110011100010",
1292 => "1001000000001100011010001",
1293 => "1001000000000110011000010",
1294 => "0001100001100100001110001",
1295 => "0001100010100100000100011",
1296 => "0100100110011101001010001",
1297 => "0100101100011100011000011",
1298 => "0000000000001100011010001",
1299 => "0001100000000110011000010",
1300 => "0110101011001100011010001",
1301 => "0110101011000110011000010",
1302 => "0000010100110000001110001",
1303 => "0100010100010000001100011",
1304 => "0110101011001100011110001",
1305 => "0110101011000110011100010",
1306 => "0010001100010100011010001",
1307 => "0010001110010100001000011",
1308 => "0110101011001100011010001",
1309 => "0110101011000110011000010",
1310 => "0010101011001100011110001",
1311 => "0100001011000110011100010",
1312 => "0011100100010110110010001",
1313 => "0011101000010110010000011",
1314 => "0011001111010100010010001",
1315 => "0011010001010100001000010",
1316 => "0111000000001100100110001",
1317 => "1000000000000100100100011",
1318 => "0010000000001100100110001",
1319 => "0011000000000100100100011",
1320 => "0101100010001000111110001",
1321 => "0101100111001000010100011",
1322 => "0000000000101000001110001",
1323 => "0000000001101000000100011",
1324 => "0110110010010100011010001",
1325 => "0110110100010100001000011",
1326 => "0001000111001100101110001",
1327 => "0010100111000110101100010",
1328 => "0101001110010100100110001",
1329 => "0101010001010100001100011",
1330 => "0100000010001000100110001",
1331 => "0101000010000100100100010",
1332 => "0111000011010100010010001",
1333 => "0111000011001010010000010",
1334 => "0011000110011000011010001",
1335 => "0011000110001100001100010",
1336 => "0110001001001100001100010",
1337 => "0100001000010000101010001",
1338 => "0110001000001000010100010",
1339 => "0100001101001000010100010",
1340 => "0011100100001001000010001",
1341 => "0011101100001000100000010",
1342 => "0100001000010010010010001",
1343 => "0100001010010010001000010",
1344 => "0010100010011100100110001",
1345 => "0010100101011100001100011",
1346 => "0001110000100110100010001",
1347 => "0001110100100110010000010",
1348 => "0000000000010100100010001",
1349 => "0010100000001010100000010",
1350 => "0010100010100001001010001",
1351 => "0010100010010001001000010",
1352 => "0000001011110000101110001",
1353 => "0100001011010000101100011",
1354 => "0001100011100100010110001",
1355 => "0001100011010010010100010",
1356 => "0000110000100100001110001",
1357 => "0000110001100100000100011",
1358 => "0010110001100100001110001",
1359 => "0010110010100100000100011",
1360 => "0000101101010010011010001",
1361 => "0000101111010010001000011",
1362 => "0000101001101110101010001",
1363 => "0000101110101110010100010",
1364 => "0001100111100100001110001",
1365 => "0001101000100100000100011",
1366 => "0011001000011000001110001",
1367 => "0011001000001100001100010",
1368 => "0011000010000111011010001",
1369 => "0011100010000011011000011",
1370 => "0111010001010100011010001",
1371 => "0111010011010100001000011",
1372 => "0000110010010100011010001",
1373 => "0000110100010100001000011",
1374 => "0101100011001100110010001",
1375 => "0110100011000100110000011",
1376 => "0101000110001000100110001",
1377 => "0110000110000100100100010",
1378 => "0101100000001100100110001",
1379 => "0110100000000100100100011",
1380 => "0011100000001100100110001",
1381 => "0100100000000100100100011",
1382 => "0110001010010010011010001",
1383 => "0111101010000110011000011",
1384 => "0001001011001100100110001",
1385 => "0010101011000110100100010",
1386 => "0111000101000111001110001",
1387 => "0111100101000011001100011",
1388 => "0011000110010010011010001",
1389 => "0011001000010010001000011",
1390 => "0111000101000111001110001",
1391 => "0111100101000011001100011",
1392 => "0000000011001100100110001",
1393 => "0000000110001100001100011",
1394 => "0010110101100100001110001",
1395 => "0010110110100100000100011",
1396 => "0000101010100100010010001",
1397 => "0011101010001100010000011",
1398 => "0110100100010000101010001",
1399 => "1000100100001000010100010",
1400 => "0110101001001000010100010",
1401 => "0011101000010010011010001",
1402 => "0101001000000110011000011",
1403 => "0110001001010010100010001",
1404 => "0111101001000110100000011",
1405 => "0000000110001010110010001",
1406 => "0000001010001010010000011",
1407 => "0011100110011100011010001",
1408 => "0111000110001110001100010",
1409 => "0011101001001110001100010",
1410 => "0011100101000111001110001",
1411 => "0100000101000011001100011",
1412 => "0100000100011111010010001",
1413 => "0110100100001011010000011",
1414 => "0000100100011111010010001",
1415 => "0011000100001011010000011",
1416 => "0110101010001100011010001",
1417 => "0110101010000110011000010",
1418 => "0010101010001100011010001",
1419 => "0100001010000110011000010",
1420 => "0111000010001100111010001",
1421 => "1000100010000110011100010",
1422 => "0111001001000110011100010",
1423 => "0010000010001100111010001",
1424 => "0010000010000110011100010",
1425 => "0011101001000110011100010",
1426 => "0110000100001100011110001",
1427 => "0110000100000110011100010",
1428 => "0100100100001100100110001",
1429 => "0101100100000100100100011",
1430 => "0101100100010000101010001",
1431 => "0101100100001000101000010",
1432 => "0010100100010000101010001",
1433 => "0100100100001000101000010",
1434 => "0100010010010100011010001",
1435 => "0100010100010100001000011",
1436 => "0000110010101010011010001",
1437 => "0000110100101010001000011",
1438 => "0100100010011000011010001",
1439 => "0100100010001100011000010",
1440 => "0001100010011000011010001",
1441 => "0100100010001100011000010",
1442 => "0110000101011000011010001",
1443 => "1001000101001100001100010",
1444 => "0110001000001100001100010",
1445 => "0100001000001100100110001",
1446 => "0100001011001100001100011",
1447 => "0001000111101000011010001",
1448 => "0001001001101000001000011",
1449 => "0000000101011000011010001",
1450 => "0000000101001100001100010",
1451 => "0011001000001100001100010",
1452 => "0111001110010000101010001",
1453 => "1001001110001000010100010",
1454 => "0111010011001000010100010",
1455 => "0001001110010000101010001",
1456 => "0001001110001000010100010",
1457 => "0011010011001000010100010",
1458 => "0001001011101000110110001",
1459 => "0001001011010100110100010",
1460 => "0011001001011000010110001",
1461 => "0110001001001100010100010",
1462 => "0010100110100000011010001",
1463 => "0110100110010000001100010",
1464 => "0010101001010000001100010",
1465 => "0000110011010010010010001",
1466 => "0000110101010010001000010",
1467 => "0011100101011000010110001",
1468 => "0101100101001000010100011",
1469 => "0001100101011100110010001",
1470 => "0001100101001110011000010",
1471 => "0101001011001110011000010",
1472 => "0100100100010010011010001",
1473 => "0110000100000110011000011",
1474 => "0001000110100110001110001",
1475 => "0001000111100110000100011",
1476 => "1001001010001100100110001",
1477 => "1001001101001100001100011",
1478 => "0001100111100100001010001",
1479 => "0001101000100100000100010",
1480 => "1010000010001001001010001",
1481 => "1011000010000100100100010",
1482 => "1010001011000100100100010",
1483 => "0001010010101000001110001",
1484 => "0001010011101000000100011",
1485 => "0000101001101100001110001",
1486 => "0000101010101100000100011",
1487 => "0000000010001001001010001",
1488 => "0000000010000100100100010",
1489 => "0001001011000100100100010",
1490 => "1001100000001001011110001",
1491 => "1001100000000101011100010",
1492 => "0000000011001101001110001",
1493 => "0001100011000111001100010",
1494 => "1001000010001100100110001",
1495 => "1010000010000100100100011",
1496 => "0000000101010100011010001",
1497 => "0000000111010100001000011",
1498 => "0011100000011000110010001",
1499 => "0110100000001100011000010",
1500 => "0011100110001100011000010",
1501 => "0000000011110000011010001",
1502 => "0000000011011000001100010",
1503 => "0110000110011000001100010",
1504 => "0101001110001000101010001",
1505 => "0101010011001000010100010",
1506 => "0100001001001000111110001",
1507 => "0100001110001000010100011",
1508 => "0010001011100010011010001",
1509 => "0010001110100010001100010",
1510 => "0001000101100100100010001",
1511 => "0001000101010010010000010",
1512 => "0101101001010010010000010",
1513 => "0011100110011100011010001",
1514 => "0111000110001110001100010",
1515 => "0011101001001110001100010",
1516 => "0001100110011100011010001",
1517 => "0001100110001110001100010",
1518 => "0101001001001110001100010",
1519 => "1000000101000111001010001",
1520 => "1000100101000011001000011",
1521 => "0010100101000111001010001",
1522 => "0011000101000011001000011",
1523 => "0101001010011100010010001",
1524 => "0101001100011100001000010",
1525 => "0010001010010010010010001",
1526 => "0010001100010010001000010",
1527 => "0001000000100100100110001",
1528 => "0001000011100100001100011",
1529 => "0011000011011000100010001",
1530 => "0101000011001000100000011",
1531 => "0000100001010000010110001",
1532 => "0010100001001000010100010",
1533 => "0110000111001110100010001",
1534 => "0110001011001110010000010",
1535 => "0000001100101100010010001",
1536 => "0000001110101100001000010",
1537 => "0111100110001000111110001",
1538 => "0111101011001000010100011",
1539 => "0010100111001110100010001",
1540 => "0010101011001110010000010",
1541 => "0100010010010010010010001",
1542 => "0100010100010010001000010",
1543 => "0000100010101100010010001",
1544 => "0000100100101100001000010",
1545 => "1000100011001101000110001",
1546 => "1001100011000101000100011",
1547 => "0100000010010001001010001",
1548 => "0100001011010000100100010",
1549 => "1000100000001100110010001",
1550 => "1010000000000110011000010",
1551 => "1000100110000110011000010",
1552 => "0011100000001100100110001",
1553 => "0100100000000100100100011",
1554 => "0111100101010010110010001",
1555 => "0111101011010010011000010",
1556 => "0001010110100100001010001",
1557 => "0001010111100100000100010",
1558 => "0101001010011000011010001",
1559 => "1000001010001100001100010",
1560 => "0101001101001100001100010",
1561 => "0000000001001000101110001",
1562 => "0001000001000100101100010",
1563 => "1010000000001000101010001",
1564 => "1010000000000100101000010",
1565 => "0000100011001101000110001",
1566 => "0001100011000101000100011",
1567 => "0111101111010010011010001",
1568 => "0111110001010010001000011",
1569 => "0000001101010000100110001",
1570 => "0000010000010000001100011",
1571 => "1000001000001100110010001",
1572 => "1000001100001100010000011",
1573 => "0001001000001100110010001",
1574 => "0001001100001100010000011",
1575 => "0101000010001000111110001",
1576 => "0101000111001000010100011",
1577 => "0000100101100110001110001",
1578 => "0000100110100110000100011",
1579 => "0101101000010010011110001",
1580 => "0111001000000110011100011",
1581 => "0001101000011000100110001",
1582 => "0001101011011000001100011",
1583 => "0001100110100100001110001",
1584 => "0001100111100100000100011",
1585 => "0101000000001000110010001",
1586 => "0101000110001000011000010",
1587 => "0001101001100100111010001",
1588 => "0001101001010010111000010",
1589 => "0000000000001000100110001",
1590 => "0001000000000100100100010",
1591 => "0110000101001001001010001",
1592 => "0110000101000101001000010",
1593 => "0100000101001001001010001",
1594 => "0101000101000101001000010",
1595 => "0101000101001100101010001",
1596 => "0110000101000100101000011",
1597 => "0100100100001000101110001",
1598 => "0101100100000100101100010",
1599 => "0010010000100100001110001",
1600 => "0010010001100100000100011",
1601 => "0000010000101000001110001",
1602 => "0000010001101000000100011",
1603 => "0100101001001100110010001",
1604 => "0100101101001100010000011",
1605 => "0100001101010000100010001",
1606 => "0100010001010000010000010",
1607 => "0110101010000110110010001",
1608 => "0110110000000110011000010",
1609 => "0010101001011100111010001",
1610 => "0010101001001110011100010",
1611 => "0110010000001110011100010",
1612 => "0000000000110000101010001",
1613 => "0110000000011000010100010",
1614 => "0000000101011000010100010",
1615 => "0000101011100100001010001",
1616 => "0000101100100100000100010",
1617 => "1001100101001010110010001",
1618 => "1001101001001010010000011",
1619 => "0000000101001010110010001",
1620 => "0000001001001010010000011",
1621 => "1000000110010001001010001",
1622 => "1010000110001000100100010",
1623 => "1000001111001000100100010",
1624 => "0000000110010001001010001",
1625 => "0000000110001000100100010",
1626 => "0010001111001000100100010",
1627 => "0110000101011000110010001",
1628 => "1001000101001100011000010",
1629 => "0110001011001100011000010",
1630 => "0011100110001100100110001",
1631 => "0100100110000100100100011",
1632 => "0100101101001100101110001",
1633 => "0101101101000100101100011",
1634 => "0000000101011000110010001",
1635 => "0000000101001100011000010",
1636 => "0011001011001100011000010",
1637 => "0000100010101110001110001",
1638 => "0000100011101110000100011",
1639 => "0000101111100110001110001",
1640 => "0000110000100110000100011",
1641 => "0110110001010110010010001",
1642 => "0110110011010110001000010",
1643 => "0000001101010000010110001",
1644 => "0010001101001000010100010",
1645 => "0110001010010100010010001",
1646 => "0110001010001010010000010",
1647 => "0010000110010010100110001",
1648 => "0010001001010010001100011",
1649 => "0111101110010010011010001",
1650 => "0111110000010010001000011",
1651 => "0000101100010010011010001",
1652 => "0000101110010010001000011",
1653 => "0001101010101000100010001",
1654 => "0110101010010100010000010",
1655 => "0001101110010100010000010",
1656 => "0001000000010011001010001",
1657 => "0010100000000111001000011",
1658 => "0110101011010010101010001",
1659 => "1000001011000110101000011",
1660 => "0000100010010000010110001",
1661 => "0010100010001000010100010",
1662 => "0001100100101010011010001",
1663 => "0101000100001110011000011",
1664 => "0011100000010100111010001",
1665 => "0011100000001010011100010",
1666 => "0110000111001010011100010",
1667 => "0110010001011000010010001",
1668 => "0110010011011000001000010",
1669 => "0000000110101110010010001",
1670 => "0000001000101110001000010",
1671 => "0110101010010000101010001",
1672 => "1000101010001000010100010",
1673 => "0110101111001000010100010",
1674 => "0000010000100100001110001",
1675 => "0000010001100100000100011",
1676 => "0111110000010010010010001",
1677 => "0111110010010010001000010",
1678 => "0000010000010010010010001",
1679 => "0000010010010010001000010",
1680 => "0110101011001100011010001",
1681 => "0110101011000110011000010",
1682 => "0010101011001100011010001",
1683 => "0100001011000110011000010",
1684 => "0000000011110000011010001",
1685 => "0110000011011000001100010",
1686 => "0000000110011000001100010",
1687 => "0001000100100100001110001",
1688 => "0001000101100100000100011",
1689 => "0000000000110000010010001",
1690 => "0110000000011000001000010",
1691 => "0000000010011000001000010",
1692 => "0000110000100100001110001",
1693 => "0000110001100100000100011",
1694 => "0111101111010010011010001",
1695 => "0111110001010010001000011",
1696 => "0000001111010010011010001",
1697 => "0000010001010010001000011",
1698 => "0011010001100100001110001",
1699 => "0011010010100100000100011",
1700 => "0100001000001100101010001",
1701 => "0101001000000100101000011",
1702 => "0101000110001100100110001",
1703 => "0110000110000100100100011",
1704 => "0100001000001010100010001",
1705 => "0100001100001010010000010",
1706 => "0110001000001100100010001",
1707 => "0110001100001100010000010",
1708 => "0011000101001100101110001",
1709 => "0100000101000100101100011",
1710 => "0110100110010000100110001",
1711 => "0110101001010000001100011",
1712 => "0000100111101010011010001",
1713 => "0000101001101010001000011",
1714 => "0111100101000110110010001",
1715 => "0111101011000110011000010",
1716 => "0011001001010110110010001",
1717 => "0011001101010110010000011",
1718 => "0110101000010100100010001",
1719 => "1001001000001010010000010",
1720 => "0110101100001010010000010",
1721 => "0010101000011000001110001",
1722 => "0101101000001100001100010",
1723 => "0011001011100100010010001",
1724 => "0110001011001100010000011",
1725 => "0000000000101101011010001",
1726 => "0000001011101100101100010",
1727 => "0101100010001100100010001",
1728 => "0101100110001100010000010",
1729 => "0100100000001100100110001",
1730 => "0101100000000100100100011",
1731 => "0101000000001100100110001",
1732 => "0110000000000100100100011",
1733 => "0100000011001100111010001",
1734 => "0100000011000110011100010",
1735 => "0101101010000110011100010",
1736 => "0001101010100100100010001",
1737 => "0100101010001100100000011",
1738 => "0101000000000110111010001",
1739 => "0101000111000110011100010",
1740 => "0010000011100001010010001",
1741 => "0010001101100000101000010",
1742 => "0100100100001100101010001",
1743 => "0101100100000100101000011",
1744 => "0010100000100000010010001",
1745 => "0010100010100000001000010",
1746 => "0001000101100100010010001",
1747 => "0100000101001100010000011",
1748 => "0110100000001100100110001",
1749 => "0111100000000100100100011",
1750 => "0100000100010000010110001",
1751 => "0110000100001000010100010",
1752 => "0110001010010100010010001",
1753 => "0110001010001010010000010",
1754 => "0001001010010100010010001",
1755 => "0011101010001010010000010",
1756 => "0011101011011000010110001",
1757 => "0101101011001000010100011",
1758 => "0001101010010000101010001",
1759 => "0001101010001000010100010",
1760 => "0011101111001000010100010",
1761 => "0101101100010010100010001",
1762 => "0111001100000110100000011",
1763 => "0000010101110000001110001",
1764 => "0100010101010000001100011",
1765 => "0001110100100100010010001",
1766 => "0100110100001100010000011",
1767 => "0000101111010010011010001",
1768 => "0000110001010010001000011",
1769 => "0101110001010100010010001",
1770 => "0101110011010100001000010",
1771 => "0100101100001000110010001",
1772 => "0100110010001000011000010",
1773 => "0100100110010010011010001",
1774 => "0110000110000110011000011",
1775 => "0000101101001100100110001",
1776 => "0000110000001100001100011",
1777 => "0011010000011000010010001",
1778 => "0011010010011000001000010",
1779 => "0000100101101000001110001",
1780 => "0000100110101000000100011",
1781 => "0100000001010010100110001",
1782 => "0100000100010010001100011",
1783 => "0001010011010010010010001",
1784 => "0001010101010010001000010",
1785 => "0101100001001001001010001",
1786 => "0101100111001000011000011",
1787 => "0011100010010000110010001",
1788 => "0011100010001000011000010",
1789 => "0101101000001000011000010",
1790 => "0101101010010010100010001",
1791 => "0111001010000110100000011",
1792 => "0010101011011000010110001",
1793 => "0100101011001000010100011",
1794 => "0101101001010010011010001",
1795 => "0111001001000110011000011",
1796 => "0010101010001100100110001",
1797 => "0011101010000100100100011",
1798 => "0010000111001010110010001",
1799 => "0010001011001010010000011",
1800 => "0001000000101010011010001",
1801 => "0100100000001110011000011",
1802 => "0011100110010100011010001",
1803 => "0011101000010100001000011",
1804 => "0100100000001100111110001",
1805 => "0101100000000100111100011",
1806 => "0001000010100100001010001",
1807 => "0001000011100100000100010",
1808 => "0100010001010000011010001",
1809 => "0100010100010000001100010",
1810 => "0001100000100100001010001",
1811 => "0001100001100100000100010",
1812 => "0100000000010010011010001",
1813 => "0101100000000110011000011",
1814 => "0000010001100100001110001",
1815 => "0000010010100100000100011",
1816 => "0011000111011000010110001",
1817 => "0101000111001000010100011",
1818 => "0000000011001100100110001",
1819 => "0001000011000100100100011",
1820 => "1010000010001000100110001",
1821 => "1010000010000100100100010",
1822 => "0000000010001000100110001",
1823 => "0001000010000100100100010",
1824 => "0000000001110000010010001",
1825 => "0110000001011000001000010",
1826 => "0000000011011000001000010",
1827 => "0000010000010010011010001",
1828 => "0000010010010010001000011",
1829 => "0111001101010010011010001",
1830 => "0111001111010010001000011",
1831 => "0000001111100110001110001",
1832 => "0000010000100110000100011",
1833 => "0000100101101100110010001",
1834 => "0110000101010110011000010",
1835 => "0000101011010110011000010",
1836 => "0010101101001100011010001",
1837 => "0100001101000110011000010",
1838 => "0010000010101000001110001",
1839 => "0010000011101000000100011",
1840 => "0100001110001100101010001",
1841 => "0101001110000100101000011",
1842 => "0011001100100000011010001",
1843 => "0111001100010000001100010",
1844 => "0011001111010000001100010",
1845 => "0001001101010000100110001",
1846 => "0001010000010000001100011",
1847 => "0101101000001100111010001",
1848 => "0111001000000110011100010",
1849 => "0101101111000110011100010",
1850 => "0001001100100000011010001",
1851 => "0001001100010000001100010",
1852 => "0101001111010000001100010",
1853 => "0010110000100000100010001",
1854 => "0010110100100000010000010",
1855 => "0100100001001000110010001",
1856 => "0100100111001000011000010",
1857 => "0100000010010000101010001",
1858 => "0110000010001000010100010",
1859 => "0100000111001000010100010",
1860 => "0011000110011000011010001",
1861 => "0011000110001100001100010",
1862 => "0110001001001100001100010",
1863 => "0101000111001100100110001",
1864 => "0110000111000100100100011",
1865 => "0000000000010000110010001",
1866 => "0000000000001000011000010",
1867 => "0010000110001000011000010",
1868 => "1001001000001100100110001",
1869 => "1001001011001100001100011",
1870 => "0001001100001100011010001",
1871 => "0010101100000110011000010",
1872 => "0001110101101010001110001",
1873 => "0101010101001110001100011",
1874 => "0001000000100000011010001",
1875 => "0001000011100000001100010",
1876 => "0110100110001110011010001",
1877 => "0110101001001110001100010",
1878 => "0011000100001000111010001",
1879 => "0011001011001000011100010",
1880 => "0100100111001100100110001",
1881 => "0101100111000100100100011",
1882 => "0011101000001100111010001",
1883 => "0011101000000110011100010",
1884 => "0101001111000110011100010",
1885 => "1001001000001001000010001",
1886 => "1001010000001000100000010",
1887 => "0100101110001100101010001",
1888 => "0101101110000100101000011",
1889 => "0011001011011000010110001",
1890 => "0101001011001000010100011",
1891 => "0000001100101110001110001",
1892 => "0000001101101110000100011",
1893 => "0110100000001100110010001",
1894 => "0111100000000100110000011",
1895 => "0000001010011000010110001",
1896 => "0010001010001000010100011",
1897 => "0110100010010100010010001",
1898 => "0110100100010100001000010",
1899 => "0010100000001100110010001",
1900 => "0011100000000100110000011",
1901 => "0101100110010010011010001",
1902 => "0111000110000110011000011",
1903 => "0010000110010010011010001",
1904 => "0011100110000110011000011",
1905 => "0011001011100100110110001",
1906 => "0110001011001100110100011",
1907 => "0000001011100100110110001",
1908 => "0011001011001100110100011",
1909 => "0110010000011000011010001",
1910 => "1000010000001000011000011",
1911 => "0000000110101010001110001",
1912 => "0000000111101010000100011",
1913 => "0110010000011000011010001",
1914 => "1000010000001000011000011",
1915 => "0010100111001100111010001",
1916 => "0010101110001100011100010",
1917 => "0010101010100110001010001",
1918 => "0010101011100110000100010",
1919 => "0010100100011100010010001",
1920 => "0010100110011100001000010",
1921 => "0001110010100100010010001",
1922 => "0100110010001100010000011",
1923 => "0011100000001000100110001",
1924 => "0100100000000100100100010",
1925 => "0110100011010110010010001",
1926 => "0110100101010110001000010",
1927 => "0001000000010010011010001",
1928 => "0010100000000110011000011",
1929 => "1001100001001001011110001",
1930 => "1001100001000101011100010",
1931 => "0000100001001001011110001",
1932 => "0001100001000101011100010",
1933 => "0010110000100100001110001",
1934 => "0010110001100100000100011",
1935 => "0000000011010110010010001",
1936 => "0000000101010110001000010",
1937 => "0001010000101000001110001",
1938 => "0001010001101000000100011",
1939 => "0010100011011010010010001",
1940 => "0010100101011010001000010",
1941 => "0000101001101100111110001",
1942 => "0000101001010110111100010",
1943 => "0001100100011100001110001",
1944 => "0101000100001110001100010",
1945 => "0100000111010100010010001",
1946 => "0100000111001010010000010",
1947 => "0011000111010100010010001",
1948 => "0101100111001010010000010",
1949 => "0101000100001100100110001",
1950 => "0110000100000100100100011",
1951 => "0000101100010010011010001",
1952 => "0010001100000110011000011",
1953 => "0100000011010000101010001",
1954 => "0110000011001000010100010",
1955 => "0100001000001000010100010",
1956 => "0001100110100000011010001",
1957 => "0001100110010000001100010",
1958 => "0101101001010000001100010",
1959 => "0010100110011100011010001",
1960 => "0010101001011100001100010",
1961 => "0010000011010010011010001",
1962 => "0010000101010010001000011",
1963 => "0011000011100100001010001",
1964 => "0011000100100100000100010",
1965 => "0011100110010010011010001",
1966 => "0101000110000110011000011",
1967 => "0000000001110000001110001",
1968 => "0000000010110000000100011",
1969 => "0000010001010100011010001",
1970 => "0000010011010100001000011",
1971 => "0001110010100100001110001",
1972 => "0001110011100100000100011",
1973 => "0001000101001101000010001",
1974 => "0001000101000110100000010",
1975 => "0010101101000110100000010",
1976 => "0011100110010110011010001",
1977 => "0011101000010110001000011",
1978 => "0010100010011001011010001",
1979 => "0010101101011000101100010",
1980 => "0101000111001000101010001",
1981 => "0101001100001000010100010",
1982 => "0100100000001001001010001",
1983 => "0100100110001000011000011",
1984 => "1001001000001100100110001",
1985 => "1001001011001100001100011",
1986 => "0010000111011110101010001",
1987 => "0100100111001010101000011",
1988 => "0101000101001100100110001",
1989 => "0110000101000100100100011",
1990 => "0100101001001100101010001",
1991 => "0101101001000100101000011",
1992 => "0101101110001100101010001",
1993 => "0110101110000100101000011",
1994 => "0011101110001100101010001",
1995 => "0100101110000100101000011",
1996 => "0010001000100000100110001",
1997 => "0010001011100000001100011",
1998 => "0001001011101000001110001",
1999 => "0001001100101000000100011",
2000 => "0110100000001000110110001",
2001 => "0110100000000100110100010",
2002 => "0011100000001000110110001",
2003 => "0100100000000100110100010",
2004 => "0001100001100100011110001",
2005 => "0100100001001100011100011",
2006 => "0000101011001100100110001",
2007 => "0000101110001100001100011",
2008 => "0100010010010010011010001",
2009 => "0100010100010010001000011",
2010 => "0001101001011110011010001",
2011 => "0001101011011110001000011",
2012 => "0010101010100110001010001",
2013 => "0010101011100110000100010",
2014 => "0100000110001111000010001",
2015 => "0100001110001110100000010",
2016 => "0100101110010010011010001",
2017 => "0100110000010010001000011",
2018 => "0000000111010000110010001",
2019 => "0000001011010000010000011",
2020 => "0011000100100100001110001",
2021 => "0011000101100100000100011",
2022 => "0000010000011000011010001",
2023 => "0010010000001000011000011",
2024 => "0110101101010010010010001",
2025 => "0110101111010010001000010",
2026 => "0010101000011100111010001",
2027 => "0010101000001110011100010",
2028 => "0110001111001110011100010",
2029 => "0000110000101100011010001",
2030 => "0110010000010110001100010",
2031 => "0000110011010110001100010",
2032 => "0100100000001100100110001",
2033 => "0101100000000100100100011",
2034 => "0100100101010100101010001",
2035 => "0111000101001010010100010",
2036 => "0100101010001010010100010",
2037 => "0010100101010100101010001",
2038 => "0010100101001010010100010",
2039 => "0101001010001010010100010",
2040 => "0010000110100000011010001",
2041 => "0110000110010000001100010",
2042 => "0010001001010000001100010",
2043 => "0000000111001100100110001",
2044 => "0000001010001100001100011",
2045 => "1000001010010000111010001",
2046 => "1010001010001000011100010",
2047 => "1000010001001000011100010",
2048 => "0100101100001100110010001",
2049 => "0100110010001100011000010",
2050 => "0100001010010000110010001",
2051 => "0110001010001000011000010",
2052 => "0100010000001000011000010",
2053 => "0100000000001000100110001",
2054 => "0101000000000100100100010",
2055 => "0101000100010001000010001",
2056 => "0111000100001000100000010",
2057 => "0101001100001000100000010",
2058 => "0011101010010100011010001",
2059 => "0011101100010100001000011",
2060 => "0010100110011100111010001",
2061 => "0110000110001110011100010",
2062 => "0010101101001110011100010",
2063 => "0001001011101000001010001",
2064 => "0001001100101000000100010",
2065 => "1001001000001001000010001",
2066 => "1001010000001000100000010",
2067 => "0000101011011000101010001",
2068 => "0000101011001100010100010",
2069 => "0011110000001100010100010",
2070 => "0011001001011000010010001",
2071 => "0011001011011000001000010",
2072 => "0100101100001100011110001",
2073 => "0110001100000110011100010",
2074 => "0101000100010001000010001",
2075 => "0111000100001000100000010",
2076 => "0101001100001000100000010",
2077 => "0011000100010001000010001",
2078 => "0011000100001000100000010",
2079 => "0101001100001000100000010",
2080 => "0100001001010010011010001",
2081 => "0101101001000110011000011",
2082 => "0000100101100000110010001",
2083 => "0000100101010000011000010",
2084 => "0100101011010000011000010",
2085 => "0100101001001100100010001",
2086 => "0100101001000110100000010",
2087 => "0011000000000111001010001",
2088 => "0011100000000011001000011",
2089 => "1000101001001010111010001",
2090 => "1000110000001010011100010",
2091 => "0001001001001010111010001",
2092 => "0001010000001010011100010",
2093 => "0011100100010100011010001",
2094 => "0011100111010100001100010",
2095 => "0000100011101111001010001",
2096 => "0000101001101110011000011",
2097 => "0000100001101010001110001",
2098 => "0100000001001110001100011",
2099 => "0100100110001100100110001",
2100 => "0101100110000100100100011",
2101 => "0001110010011000011010001",
2102 => "0001110010001100001100010",
2103 => "0100110101001100001100010",
2104 => "1000001000010001000010001",
2105 => "1010001000001000100000010",
2106 => "1000010000001000100000010",
2107 => "0000010011110000010010001",
2108 => "0100010011010000010000011",
2109 => "1000001000010001000010001",
2110 => "1010001000001000100000010",
2111 => "1000010000001000100000010",
2112 => "0000001000010001000010001",
2113 => "0000001000001000100000010",
2114 => "0010010000001000100000010",
2115 => "0100001100010000101010001",
2116 => "0100010001010000010100010",
2117 => "0010100111001010100010001",
2118 => "0010101011001010010000010",
2119 => "0010000001100110001010001",
2120 => "0010000010100110000100010",
2121 => "0000001100110000100110001",
2122 => "0100001100010000100100011",
2123 => "0011000000011010100010001",
2124 => "0011000100011010010000010",
2125 => "0000000000110000001110001",
2126 => "0000000001110000000100011",
2127 => "1010000011001000101110001",
2128 => "1010000011000100101100010",
2129 => "0100000110001100100110001",
2130 => "0101000110000100100100011",
2131 => "0011001011011000100010001",
2132 => "0110001011001100010000010",
2133 => "0011001111001100010000010",
2134 => "0000001000011000011010001",
2135 => "0000001000001100001100010",
2136 => "0011001011001100001100010",
2137 => "0011010001100100001110001",
2138 => "0011010010100100000100011",
2139 => "0000001110010010011010001",
2140 => "0000010000010010001000011",
2141 => "1010000011001000100110001",
2142 => "1010000011000100100100010",
2143 => "0000000011001000100110001",
2144 => "0001000011000100100100010",
2145 => "0111100000010011001110001",
2146 => "1001000000000111001100011",
2147 => "0000000000010011001110001",
2148 => "0001100000000111001100011",
2149 => "0110101011001100100010001",
2150 => "0110101011000110100000010",
2151 => "0010101011001100100010001",
2152 => "0100001011000110100000010",
2153 => "0010101011100110001110001",
2154 => "0010101100100110000100011",
2155 => "0001110100100100010010001",
2156 => "0100110100001100010000011",
2157 => "0011000110100000011010001",
2158 => "0011001000100000001000011",
2159 => "0011000000010010011010001",
2160 => "0100100000000110011000011",
2161 => "0101000011001000111010001",
2162 => "0101001010001000011100010",
2163 => "0000100101011110110010001",
2164 => "0000101011011110011000010",
2165 => "0101101100010000010110001",
2166 => "0101101100001000010100010",
2167 => "0010100000001100100110001",
2168 => "0011100000000100100100011",
2169 => "0110000000001100100110001",
2170 => "0111000000000100100100011",
2171 => "0010100101011000100010001",
2172 => "0010100101001100010000010",
2173 => "0101101001001100010000010",
2174 => "0110101100010110011010001",
2175 => "0110101110010110001000011",
2176 => "0000001101101010001110001",
2177 => "0000001110101010000100011",
2178 => "0100000001010000110010001",
2179 => "0110000001001000011000010",
2180 => "0100000111001000011000010",
2181 => "0000100000001100110010001",
2182 => "0000100000000110011000010",
2183 => "0010000110000110011000010",
2184 => "0001000010101010001010001",
2185 => "0001000011101010000100010",
2186 => "0001000010100110001110001",
2187 => "0001000011100110000100011",
2188 => "1000101010001100111010001",
2189 => "1010001010000110011100010",
2190 => "1000110001000110011100010",
2191 => "0000101010001100111010001",
2192 => "0000101010000110011100010",
2193 => "0010010001000110011100010",
2194 => "0011100110011100111010001",
2195 => "0111000110001110011100010",
2196 => "0011101101001110011100010",
2197 => "0000001100010010011010001",
2198 => "0000001110010010001000011",
2199 => "0111101110010000100110001",
2200 => "0111110001010000001100011",
2201 => "0000100001101100010010001",
2202 => "0000100001010110001000010",
2203 => "0110000011010110001000010",
2204 => "0100101011010010011010001",
2205 => "0100101101010010001000011",
2206 => "0000001111100100001110001",
2207 => "0000010000100100000100011",
2208 => "1000001110001110100110001",
2209 => "1000010001001110001100011",
2210 => "0010000011100000010010001",
2211 => "0110000011010000010000010",
2212 => "0011100110011000010110001",
2213 => "0011100110001100010100010",
2214 => "0100100110001000100110001",
2215 => "0101100110000100100100010",
2216 => "0110000001001000101010001",
2217 => "0110000001000100101000010",
2218 => "0100000001001000101010001",
2219 => "0101000001000100101000010",
2220 => "0111101111001100100110001",
2221 => "0111110010001100001100011",
2222 => "0001101111001100100110001",
2223 => "0001110010001100001100011",
2224 => "0111100001000111001110001",
2225 => "1000000001000011001100011",
2226 => "0000100011001100100110001",
2227 => "0001100011000100100100011",
2228 => "0111100000000111001110001",
2229 => "1000000000000011001100011",
2230 => "0011000011011000010010001",
2231 => "0110000011001100010000010",
2232 => "0101000101001000100110001",
2233 => "0101000101000100100100010",
2234 => "0011000000000111001110001",
2235 => "0011100000000011001100011",
2236 => "0101100001000110110010001",
2237 => "0101100111000110011000010",
2238 => "0011000111010100010110001",
2239 => "0101100111001010010100010",
2240 => "0101100011000111001010001",
2241 => "0110000011000011001000011",
2242 => "0100100011001100110010001",
2243 => "0101100011000100110000011",
2244 => "0001100111100110001110001",
2245 => "0001101000100110000100011",
2246 => "0001000111100100001110001",
2247 => "0001001000100100000100011",
2248 => "0001101101100100010010001",
2249 => "0110001101010010001000010",
2250 => "0001101111010010001000010",
2251 => "0001100101001100100110001",
2252 => "0010100101000100100100011",
2253 => "0010000001101000010010001",
2254 => "0111000001010100001000010",
2255 => "0010000011010100001000010",
2256 => "0000000001101000010010001",
2257 => "0000000001010100001000010",
2258 => "0101000011010100001000010",
2259 => "0101001111001100011010001",
2260 => "0101001111000110011000010",
2261 => "0000000010110000100010001",
2262 => "0100000010010000100000011",
2263 => "0010100101100100001110001",
2264 => "0010100110100100000100011",
2265 => "0100001111001100011010001",
2266 => "0101101111000110011000010",
2267 => "0101101100010000010110001",
2268 => "0101101100001000010100010",
2269 => "0010101100010000010110001",
2270 => "0100101100001000010100010",
2271 => "0010100000011100011010001",
2272 => "0010100010011100001000011",
2273 => "0101000010001000111110001",
2274 => "0101000111001000010100011",
2275 => "0101000111001010110010001",
2276 => "0101001011001010010000011",
2277 => "0011101001010000111010001",
2278 => "0011101001001000011100010",
2279 => "0101110000001000011100010",
2280 => "0000100101101100011010001",
2281 => "0110000101010110001100010",
2282 => "0000101000010110001100010",
2283 => "0000000101001100011010001",
2284 => "0000001000001100001100010",
2285 => "0110010001010010010010001",
2286 => "0110010011010010001000010",
2287 => "0001010010100110001110001",
2288 => "0001010011100110000100011",
2289 => "0110010001010010010010001",
2290 => "0110010011010010001000010",
2291 => "0000110001100100001110001",
2292 => "0000110010100100000100011",
2293 => "0110010001010010010010001",
2294 => "0110010011010010001000010",
2295 => "0000000000110000001110001",
2296 => "0000000001110000000100011",
2297 => "0010100000011100010010001",
2298 => "0010100010011100001000010",
2299 => "0011001110010010011010001",
2300 => "0011010000010010001000011",
2301 => "0111001101001100100110001",
2302 => "0111010000001100001100011",
2303 => "0010110100011010010010001",
2304 => "0010110110011010001000010",
2305 => "0100101001001100110010001",
2306 => "0100101101001100010000011",
2307 => "0000101010101010001110001",
2308 => "0100001010001110001100011",
2309 => "0100001000010010011010001",
2310 => "0101101000000110011000011",
2311 => "0001101010010010011110001",
2312 => "0011001010000110011100011",
2313 => "0110001010010100100010001",
2314 => "1000101010001010010000010",
2315 => "0110001110001010010000010",
2316 => "0000001111110000001110001",
2317 => "0100001111010000001100011",
2318 => "0100000101010010011010001",
2319 => "0100000111010010001000011",
2320 => "0010001101001100100110001",
2321 => "0010010000001100001100011",
2322 => "0110010001010010010010001",
2323 => "0110010011010010001000010",
2324 => "0100101100001100011010001",
2325 => "0100101111001100001100010",
2326 => "0100101001011100101010001",
2327 => "1000001001001110010100010",
2328 => "0100101110001110010100010",
2329 => "0000101001011100101010001",
2330 => "0000101001001110010100010",
2331 => "0100001110001110010100010",
2332 => "0100000111010011000110001",
2333 => "0101100111000111000100011",
2334 => "0001100100001101010010001",
2335 => "0001100100000110101000010",
2336 => "0011001110000110101000010",
2337 => "0011101000010100010010001",
2338 => "0011101000001010010000010",
2339 => "0101000111001000100110001",
2340 => "0110000111000100100100010",
2341 => "0101001111001100100110001",
2342 => "0110001111000100100100011",
2343 => "0001101000001101000010001",
2344 => "0001101000000110100000010",
2345 => "0011010000000110100000010",
2346 => "0110010001010010010010001",
2347 => "0110010011010010001000010",
2348 => "0001110001010010010010001",
2349 => "0001110011010010001000010",
2350 => "0101000001010010011010001",
2351 => "0110100001000110011000011",
2352 => "0010100111001000101010001",
2353 => "0010101100001000010100010",
2354 => "0011100101011000011010001",
2355 => "0101100101001000011000011",
2356 => "0011000100010010100010001",
2357 => "0100100100000110100000011",
2358 => "0110010000010100100010001",
2359 => "1000110000001010010000010",
2360 => "0110010100001010010000010",
2361 => "0001010000010100100010001",
2362 => "0001010000001010010000010",
2363 => "0011110100001010010000010",
2364 => "0000000000110000010010001",
2365 => "0110000000011000001000010",
2366 => "0000000010011000001000010",
2367 => "0000000110010010011010001",
2368 => "0000001000010010001000011",
2369 => "0000000100110000011010001",
2370 => "0110000100011000001100010",
2371 => "0000000111011000001100010",
2372 => "0010100000010110010010001",
2373 => "0010100010010110001000010",
2374 => "0000100001101100010010001",
2375 => "0110000001010110001000010",
2376 => "0000100011010110001000010",
2377 => "0100100110001101001010001",
2378 => "0100101111001100100100010",
2379 => "0001001001101000010010001",
2380 => "0001001011101000001000010",
2381 => "0010100010011100111010001",
2382 => "0010101001011100011100010",
2383 => "0010000010100000011010001",
2384 => "0010000101100000001100010",
2385 => "0001000011100110001110001",
2386 => "0001000100100110000100011",
2387 => "0011100001010100010010001",
2388 => "0011100011010100001000010",
2389 => "0000001001001000111110001",
2390 => "0000001110001000010100011",
2391 => "0001001010101010001110001",
2392 => "0001001011101010000100011",
2393 => "0001100000001100011010001",
2394 => "0011000000000110011000010",
2395 => "0011000100011100100110001",
2396 => "0011000111011100001100011",
2397 => "0100100001001100100110001",
2398 => "0101100001000100100100011",
2399 => "0111101000010010100110001",
2400 => "0111101011010010001100011",
2401 => "0100000000001001010110001",
2402 => "0100000111001000011100011",
2403 => "0001110110100110001010001",
2404 => "0001110111100110000100010",
2405 => "0001001111101000001110001",
2406 => "0001010000101000000100011",
2407 => "1001100000001000110110001",
2408 => "1001100000000100110100010",
2409 => "0000100111010000100010001",
2410 => "0000101011010000010000010",
2411 => "0111001110001100100110001",
2412 => "0111010001001100001100011",
2413 => "0010001110001100100110001",
2414 => "0010010001001100001100011",
2415 => "0111000101001000101010001",
2416 => "0111000101000100101000010",
2417 => "0011000101001000101010001",
2418 => "0100000101000100101000010",
2419 => "0111000101001100011010001",
2420 => "0111001000001100001100010",
2421 => "0010000101001100011010001",
2422 => "0010001000001100001100010",
2423 => "0000000010110001010110001",
2424 => "0100000010010001010100011",
2425 => "0000100010001100110110001",
2426 => "0001100010000100110100011",
2427 => "1010000000001001010110001",
2428 => "1010000000000101010100010",
2429 => "0000000100001001010010001",
2430 => "0001000100000101010000010",
2431 => "0100010000010010011010001",
2432 => "0100010010010010001000011",
2433 => "0011100000001100100110001",
2434 => "0100100000000100100100011",
2435 => "1000001100001110100110001",
2436 => "1000001111001110001100011",
2437 => "0010110101011100001110001",
2438 => "0110010101001110001100010",
2439 => "0101100101001100100110001",
2440 => "0101100101000110100100010",
2441 => "0101000101001000101010001",
2442 => "0110000101000100101000010",
2443 => "0101000110001100100110001",
2444 => "0110000110000100100100011",
2445 => "0011100101001100100110001",
2446 => "0101000101000110100100010",
2447 => "0111001110010100010010001",
2448 => "0111010000010100001000010",
2449 => "0010100101011100111010001",
2450 => "0010100101001110011100010",
2451 => "0110001100001110011100010",
2452 => "0110001000011000011010001",
2453 => "1001001000001100001100010",
2454 => "0110001011001100001100010",
2455 => "0011000110011000110010001",
2456 => "0011000110001100011000010",
2457 => "0110001100001100011000010",
2458 => "0101101101001100101010001",
2459 => "0110101101000100101000011",
2460 => "0000101010101000100010001",
2461 => "0000101010010100010000010",
2462 => "0101101110010100010000010",
2463 => "0111101101010010011010001",
2464 => "0111101111010010001000011",
2465 => "0100100000001100100110001",
2466 => "0100100011001100001100011",
2467 => "0101000001001010111010001",
2468 => "0101001000001010011100010",
2469 => "0001100100100000011010001",
2470 => "0001100110100000001000011",
2471 => "1000000011010000100110001",
2472 => "1000000110010000001100011",
2473 => "0011101101001100101010001",
2474 => "0100101101000100101000011",
2475 => "0111101101010010011010001",
2476 => "0111101111010010001000011",
2477 => "0000001101010010011010001",
2478 => "0000001111010010001000011",
2479 => "0110110000010010011010001",
2480 => "0110110010010010001000011",
2481 => "0001010000010010011010001",
2482 => "0001010010010010001000011",
2483 => "0010110000100100001110001",
2484 => "0010110001100100000100011",
2485 => "0000110000100100001110001",
2486 => "0000110001100100000100011",
2487 => "0010100000100100001110001",
2488 => "0010100001100100000100011",
2489 => "0000100001100110001010001",
2490 => "0000100010100110000100010",
2491 => "0111000010001100101110001",
2492 => "1000000010000100101100011",
2493 => "0010001111011110011010001",
2494 => "0100101111001010011000011",
2495 => "0111000010001100101110001",
2496 => "1000000010000100101100011",
2497 => "0010000010001100101110001",
2498 => "0011000010000100101100011",
2499 => "1001000010001100100110001",
2500 => "1001000101001100001100011",
2501 => "0000100010101100010010001",
2502 => "0000100010010110001000010",
2503 => "0110000100010110001000010",
2504 => "0001000000101010110010001",
2505 => "0100100000001110110000011",
2506 => "0000001100100100001110001",
2507 => "0000001101100100000100011",
2508 => "0110000010001100100110001",
2509 => "0111000010000100100100011",
2510 => "0001101010100100001110001",
2511 => "0001101011100100000100011",
2512 => "1000000011010000100110001",
2513 => "1000000110010000001100011",
2514 => "0001100111100100001110001",
2515 => "0001101000100100000100011",
2516 => "0100101011001100100110001",
2517 => "0101101011000100100100011",
2518 => "0100101000001100100110001",
2519 => "0101101000000100100100011",
2520 => "0111100000000101001010001",
2521 => "0111100000000011001000010",
2522 => "0011100000000101001010001",
2523 => "0100000000000011001000010",
2524 => "1000100011001110100110001",
2525 => "1000100110001110001100011",
2526 => "0001110010010010011010001",
2527 => "0001110100010010001000011",
2528 => "0001110010101010001110001",
2529 => "0001110011101010000100011",
2530 => "0000000011001110100110001",
2531 => "0000000110001110001100011",
2532 => "0001000111101100001110001",
2533 => "0001001000101100000100011",
2534 => "0000000011110001000010001",
2535 => "0000000011011000100000010",
2536 => "0110001011011000100000010",
2537 => "0110110001010010010010001",
2538 => "0110110011010010001000010",
2539 => "0010100101011000100010001",
2540 => "0010100101001100010000010",
2541 => "0101101001001100010000010",
2542 => "0010100110011100011010001",
2543 => "0110000110001110001100010",
2544 => "0010101001001110001100010",
2545 => "0010110000011100011010001",
2546 => "0010110000001110001100010",
2547 => "0110010011001110001100010",
2548 => "1001000010001100100110001",
2549 => "1001000101001100001100011",
2550 => "0000000010001100100110001",
2551 => "0000000101001100001100011",
2552 => "0001100100101000101010001",
2553 => "0110100100010100010100010",
2554 => "0001101001010100010100010",
2555 => "0001001101010010100010001",
2556 => "0010101101000110100000011",
2557 => "0001000001101010111110001",
2558 => "0100100001001110111100011",
2559 => "0010101100011100100010001",
2560 => "0110001100001110100000010",
2561 => "0011000111011000010010001",
2562 => "0011000111001100010000010",
2563 => "0011000101010010011010001",
2564 => "0100100101000110011000011",
2565 => "0110101011001100011010001",
2566 => "0110101011000110011000010",
2567 => "0010101011001100011010001",
2568 => "0100001011000110011000010",
2569 => "0011000100100100001010001",
2570 => "0011000101100100000100010",
2571 => "0000000010001100101110001",
2572 => "0001000010000100101100011",
2573 => "1001000000001100111110001",
2574 => "1010000000000100111100011",
2575 => "0000000000001100110110001",
2576 => "0001000000000100110100011",
2577 => "0110000000001100100110001",
2578 => "0111000000000100100100011",
2579 => "0011000000001100100110001",
2580 => "0100000000000100100100011",
2581 => "0000000010110000010010001",
2582 => "0100000010010000010000011",
2583 => "0001101101100100010010001",
2584 => "0110001101010010010000010",
2585 => "0100100111010100010010001",
2586 => "0100100111001010010000010",
2587 => "0010101000011000001110001",
2588 => "0101101000001100001100010",
2589 => "0010001110100110001110001",
2590 => "0010001111100110000100011",
2591 => "0101000000001001010010001",
2592 => "0101001010001000101000010",
2593 => "0100001111010010011010001",
2594 => "0100010001010010001000011",
2595 => "0001001001011110010010001",
2596 => "0011101001001010010000011",
2597 => "0100000100011000011110001",
2598 => "0110000100001000011100011",
2599 => "0000001010001100100110001",
2600 => "0000001101001100001100011",
2601 => "1001000101001100100110001",
2602 => "1001001000001100001100011",
2603 => "0000010010100000011010001",
2604 => "0000010010010000001100010",
2605 => "0100010101010000001100010",
2606 => "0100110010011100011010001",
2607 => "1000010010001110001100010",
2608 => "0100110101001110001100010",
2609 => "0000110100101000010010001",
2610 => "0000110100010100001000010",
2611 => "0101110110010100001000010",
2612 => "0001001000101000011010001",
2613 => "0110001000010100001100010",
2614 => "0001001011010100001100010",
2615 => "0011101000001100100110001",
2616 => "0100101000000100100100011",
2617 => "0100000101011000100010001",
2618 => "0110000101001000100000011",
2619 => "0010000101011000100010001",
2620 => "0100000101001000100000011",
2621 => "0101000110001100100110001",
2622 => "0110000110000100100100011",
2623 => "0001000000001101000010001",
2624 => "0010000000000101000000011",
2625 => "0111100100001100110010001",
2626 => "0111101000001100010000011",
2627 => "0001100100001100110010001",
2628 => "0001101000001100010000011",
2629 => "0111101100010010011010001",
2630 => "0111101110010010001000011",
2631 => "0010000000011111011010001",
2632 => "0010001011011110101100010",
2633 => "0111101100010010011010001",
2634 => "0111101110010010001000011",
2635 => "0000001100010010011010001",
2636 => "0000001110010010001000011",
2637 => "0111101111010010011010001",
2638 => "0111110001010010001000011",
2639 => "0000001111010010011010001",
2640 => "0000010001010010001000011",
2641 => "0101000000010000101010001",
2642 => "0111000000001000010100010",
2643 => "0101000101001000010100010",
2644 => "0000100000001001000010001",
2645 => "0001100000000101000000010",
2646 => "0011100110010100011010001",
2647 => "0011101000010100001000011",
2648 => "0101001100001000101010001",
2649 => "0101010001001000010100010",
2650 => "0100000100010100011010001",
2651 => "0100000110010100001000011",
2652 => "0001110110100100001010001",
2653 => "0110010110010010001000010",
2654 => "0011100111010110011010001",
2655 => "0011101001010110001000011",
2656 => "0000000000011000101010001",
2657 => "0000000000001100010100010",
2658 => "0011000101001100010100010",
2659 => "0101000001011000011010001",
2660 => "1000000001001100001100010",
2661 => "0101000100001100001100010",
2662 => "0011110000010010010010001",
2663 => "0011110010010010001000010",
2664 => "0010100111011111000010001",
2665 => "0101000111001011000000011",
2666 => "0010101010011000110110001",
2667 => "0101101010001100110100010",
2668 => "0011000010011000011010001",
2669 => "0110000010001100001100010",
2670 => "0011000101001100001100010",
2671 => "0001101001011000100110001",
2672 => "0001101100011000001100011",
2673 => "1000000010010000011010001",
2674 => "1000000101010000001100010",
2675 => "0000000010010000011010001",
2676 => "0000000101010000001100010",
2677 => "0000000011110000101110001",
2678 => "0000000011011000101100010",
2679 => "0000001101010000101010001",
2680 => "0000001101001000010100010",
2681 => "0010010010001000010100010",
2682 => "0101001110001000101010001",
2683 => "0101010011001000010100010",
2684 => "0101000010001001010110001",
2685 => "0101001001001000011100011",
2686 => "0010000100011110100110001",
2687 => "0010000111011110001100011",
2688 => "0000000001110000011010001",
2689 => "0100000001010000011000011",
2690 => "0100100110001011000010001",
2691 => "0100101110001010100000010",
2692 => "0001110101100100001110001",
2693 => "0100110101001100001100011",
2694 => "0011000101000110110010001",
2695 => "0011001011000110011000010",
2696 => "0101100110001000100110001",
2697 => "0101100110000100100100010",
2698 => "0010100110010010100010001",
2699 => "0100000110000110100000011",
2700 => "0010000011101000001010001",
2701 => "0010000100101000000100010",
2702 => "0001001010100100001110001",
2703 => "0100001010001100001100011",
2704 => "0011101111010100011010001",
2705 => "0011110001010100001000011",
2706 => "0000100100001001001010001",
2707 => "0000100100000100100100010",
2708 => "0001101101000100100100010",
2709 => "0110100000001100100110001",
2710 => "0111100000000100100100011",
2711 => "0010100000001100100110001",
2712 => "0011100000000100100100011",
2713 => "0101100000001100100110001",
2714 => "0110100000000100100100011",
2715 => "0011000111010010011010001",
2716 => "0100100111000110011000011",
2717 => "0001100000100100001010001",
2718 => "0001100001100100000100010",
2719 => "0000001010101000010010001",
2720 => "0000001010010100001000010",
2721 => "0101001100010100001000010",
2722 => "0101000010001000110010001",
2723 => "0101001000001000011000010",
2724 => "0011000101001100110010001",
2725 => "0011000101000110011000010",
2726 => "0100101011000110011000010",
2727 => "0011000000100101011010001",
2728 => "0111100000010010101100010",
2729 => "0011001011010010101100010",
2730 => "0000000000100101011010001",
2731 => "0000000000010010101100010",
2732 => "0100101011010010101100010",
2733 => "1001000010001100101110001",
2734 => "1010000010000100101100011",
2735 => "0000000010001100101110001",
2736 => "0001000010000100101100011",
2737 => "0101100000001100100110001",
2738 => "0110100000000100100100011",
2739 => "0000000000101000001110001",
2740 => "0000000001101000000100011",
2741 => "0001000010101000001010001",
2742 => "0001000011101000000100010",
2743 => "0000101010100100001010001",
2744 => "0000101011100100000100010",
2745 => "1001000111001100100110001",
2746 => "1001001010001100001100011",
2747 => "0000000000101100100110001",
2748 => "0000000011101100001100011",
2749 => "1000100011001100100110001",
2750 => "1000100110001100001100011",
2751 => "0000000111001100100110001",
2752 => "0000001010001100001100011",
2753 => "0000000110110000011010001",
2754 => "0000001000110000001000011",
2755 => "0000000010001100101010001",
2756 => "0001000010000100101000011",
2757 => "0101000110001100100110001",
2758 => "0110000110000100100100011",
2759 => "0011100000001100100110001",
2760 => "0100100000000100100100011",
2761 => "0111100000001100100110001",
2762 => "1000100000000100100100011",
2763 => "0001100000001100100110001",
2764 => "0010100000000100100100011",
2765 => "0111110001010010011010001",
2766 => "0111110011010010001000011",
2767 => "0000010001100100001110001",
2768 => "0000010010100100000100011",
2769 => "0111101110010010011010001",
2770 => "0111110000010010001000011",
2771 => "0000001111101110011010001",
2772 => "0000010001101110001000011",
2773 => "0010101111100100001110001",
2774 => "0010110000100100000100011",
2775 => "0000001110010010011010001",
2776 => "0000010000010010001000011",
2777 => "0100101000010000101010001",
2778 => "0110101000001000010100010",
2779 => "0100101101001000010100010",
2780 => "0001100111011110011010001",
2781 => "0100000111001010011000011",
2782 => "0100101000010000101010001",
2783 => "0110101000001000010100010",
2784 => "0100101101001000010100010",
2785 => "0010100000001100110010001",
2786 => "0100000000000110110000010",
2787 => "0100101000010000101010001",
2788 => "0110101000001000010100010",
2789 => "0100101101001000010100010",
2790 => "0100000101001100100110001",
2791 => "0101000101000100100100011",
2792 => "0101000110001001001010001",
2793 => "0110000110000100100100010",
2794 => "0101001111000100100100010",
2795 => "0010100111011000010010001",
2796 => "0101100111001100010000010",
2797 => "0100101000010000101010001",
2798 => "0110101000001000010100010",
2799 => "0100101101001000010100010",
2800 => "0011101000010000101010001",
2801 => "0011101000001000010100010",
2802 => "0101101101001000010100010",
2803 => "0101101010001100111010001",
2804 => "0111001010000110011100010",
2805 => "0101110001000110011100010",
2806 => "0100100101001101001110001",
2807 => "0110000101000111001100010",
2808 => "0011001100011000011010001",
2809 => "0110001100001100001100010",
2810 => "0011001111001100001100010",
2811 => "0000101001100100011010001",
2812 => "0000101001010010001100010",
2813 => "0101001100010010001100010",
2814 => "1000001110010000101010001",
2815 => "1010001110001000010100010",
2816 => "1000010011001000010100010",
2817 => "0000001001101100100010001",
2818 => "0000001001010110010000010",
2819 => "0101101101010110010000010",
2820 => "0100010010011000011010001",
2821 => "0111010010001100001100010",
2822 => "0100010101001100001100010",
2823 => "0000000110101001001010001",
2824 => "0000000110010100100100010",
2825 => "0101001111010100100100010",
2826 => "0001100110101000110010001",
2827 => "0110100110010100011000010",
2828 => "0001101100010100011000010",
2829 => "0000010000010100100010001",
2830 => "0000010000001010010000010",
2831 => "0010110100001010010000010",
2832 => "0011010000100100001110001",
2833 => "0011010001100100000100011",
2834 => "0000001011100110001110001",
2835 => "0000001100100110000100011",
2836 => "0111000110001100100110001",
2837 => "0111001001001100001100011",
2838 => "0000100111101100010010001",
2839 => "0000100111010110001000010",
2840 => "0110001001010110001000010",
2841 => "0110100110001110110010001",
2842 => "0110101010001110010000011",
2843 => "0010000111010110100110001",
2844 => "0010001010010110001100011",
2845 => "0110001010010100100010001",
2846 => "1000101010001010010000010",
2847 => "0110001110001010010000010",
2848 => "0001001100010010011110001",
2849 => "0010101100000110011100011",
2850 => "1000001110001100100110001",
2851 => "1000010001001100001100011",
2852 => "0001101100001100110010001",
2853 => "0001110000001100010000011",
2854 => "0111001101001100011010001",
2855 => "0111010000001100001100010",
2856 => "0100000000001100100110001",
2857 => "0101000000000100100100011",
2858 => "0100100001001101011110001",
2859 => "0101100001000101011100011",
2860 => "0000010000010010011010001",
2861 => "0000010010010010001000011",
2862 => "0010010001100100001110001",
2863 => "0010010010100100000100011",
2864 => "0010100010011010111010001",
2865 => "0010101001011010011100010",
2866 => "0111100000010000110010001",
2867 => "1001100000001000011000010",
2868 => "0111100110001000011000010",
2869 => "0000000000010000110010001",
2870 => "0000000000001000011000010",
2871 => "0010000110001000011000010",
2872 => "0100000010010000011110001",
2873 => "0100000010001000011100010",
2874 => "0000100001001100100110001",
2875 => "0001100001000100100100011",
2876 => "0111001000001100110010001",
2877 => "1000101000000110011000010",
2878 => "0111001110000110011000010",
2879 => "0010001000001100110010001",
2880 => "0010001000000110011000010",
2881 => "0011101110000110011000010",
2882 => "1000000101001010111110001",
2883 => "1000001010001010010100011",
2884 => "0001100101001010111110001",
2885 => "0001101010001010010100011",
2886 => "1001000100001100100110001",
2887 => "1001000111001100001100011",
2888 => "0000100111001100111110001",
2889 => "0000101100001100010100011",
2890 => "0101101111011000100010001",
2891 => "1000101111001100010000010",
2892 => "0101110011001100010000010",
2893 => "0000000010110000010010001",
2894 => "0000000010011000001000010",
2895 => "0110000100011000001000010",
2896 => "0111100001000101001110001",
2897 => "0111100001000011001100010",
2898 => "0011100001000101001110001",
2899 => "0100000001000011001100010",
2900 => "1011000001000101010010001",
2901 => "1011000001000011010000010",
2902 => "0000000001000101010010001",
2903 => "0000100001000011010000010",
2904 => "1001001011001100110010001",
2905 => "1010001011000100110000011",
2906 => "0000001011001100110010001",
2907 => "0001001011000100110000011",
2908 => "0001100110100100111010001",
2909 => "0001101101100100011100010",
2910 => "0011001010001110100010001",
2911 => "0011001110001110010000010",
2912 => "0011101001011000110010001",
2913 => "0011101101011000010000011",
2914 => "0001010010100100010110001",
2915 => "0101110010010010010100010",
2916 => "0010010101101000001110001",
2917 => "0010010110101000000100011",
2918 => "0100101100001100110010001",
2919 => "0100101100000110011000010",
2920 => "0110010010000110011000010",
2921 => "0010000110100100001110001",
2922 => "0010000111100100000100011",
2923 => "0001100110100100001110001",
2924 => "0001100111100100000100011",
2925 => "1001000100001100100110001",
2926 => "1001000111001100001100011",
2927 => "0001001100010010011010001",
2928 => "0001001110010010001000011",
2929 => "0010001110100100010010001",
2930 => "0110101110010010001000010",
2931 => "0010010000010010001000010",
2932 => "0011100111001100111010001",
2933 => "0011100111000110011100010",
2934 => "0101001110000110011100010",
2935 => "0011101101011000011010001",
2936 => "0110101101001100001100010",
2937 => "0011110000001100001100010",
2938 => "0011000111011000100110001",
2939 => "0101000111001000100100011",
2940 => "0110001100001100011010001",
2941 => "0110001100000110011000010",
2942 => "0000000010001000101010001",
2943 => "0000000111001000010100010",
2944 => "0100000000010010011010001",
2945 => "0101100000000110011000011",
2946 => "0001001001011000011010001",
2947 => "0001001100011000001100010",
2948 => "0110101010001100100110001",
2949 => "0110101101001100001100011",
2950 => "0010101010001100100110001",
2951 => "0010101101001100001100011",
2952 => "0100101111010010011010001",
2953 => "0100110001010010001000011",
2954 => "0010110000011000011010001",
2955 => "0010110011011000001100010",
2956 => "0001100010101000001110001",
2957 => "0001100011101000000100011",
2958 => "0001000101011000011010001",
2959 => "0011000101001000011000011",
2960 => "0101100000000111100010001",
2961 => "0110000000000011100000011",
2962 => "0001110000011110010010001",
2963 => "0100010000001010010000011",
2964 => "0100101100001100110010001",
2965 => "0100110010001100011000010",
2966 => "0000101111011000100010001",
2967 => "0000101111001100010000010",
2968 => "0011110011001100010000010",
2969 => "0111101010010000111010001",
2970 => "1001101010001000011100010",
2971 => "0111110001001000011100010",
2972 => "0000101001010000111010001",
2973 => "0000101001001000011100010",
2974 => "0010110000001000011100010",
2975 => "0100101011010010101010001",
2976 => "0100110000010010010100010",
2977 => "0011000111011000011010001",
2978 => "0011001001011000001000011",
2979 => "0101001111001100100110001",
2980 => "0110001111000100100100011",
2981 => "0011101000010010011110001",
2982 => "0101001000000110011100011",
2983 => "0101000100010000101010001",
2984 => "0111000100001000010100010",
2985 => "0101001001001000010100010",
2986 => "0010000110001100100110001",
2987 => "0010001001001100001100011",
2988 => "0000000110110000110010001",
2989 => "0100000110010000110000011",
2990 => "0001100111001100111010001",
2991 => "0011000111000110111000010",
2992 => "1001101000001010100010001",
2993 => "1001101100001010010000010",
2994 => "0000001000001010100010001",
2995 => "0000001100001010010000010",
2996 => "1000100011001100011010001",
2997 => "1000100110001100001100010",
2998 => "0000100011001100011010001",
2999 => "0000100110001100001100010",
3000 => "1001000010001100100110001",
3001 => "1001000101001100001100011",
3002 => "0000000010001100100110001",
3003 => "0000000101001100001100011",
3004 => "0001100011100100011010001",
3005 => "0001100101100100001000011",
3006 => "0001000011010010011010001",
3007 => "0001000101010010001000011",
3008 => "0100100011010100100010001",
3009 => "0111000011001010010000010",
3010 => "0100100111001010010000010",
3011 => "0010100011010100100010001",
3012 => "0010100011001010010000010",
3013 => "0101000111001010010000010",
3014 => "0101001011001100110010001",
3015 => "0101001011000110110000010",
3016 => "0100001011001100101110001",
3017 => "0101101011000110101100010",
3018 => "0011101000010100010010001",
3019 => "0011101000001010010000010",
3020 => "0100100110001100011110001",
3021 => "0110000110000110011100010",
3022 => "0010110010100100001110001",
3023 => "0010110011100100000100011",
3024 => "0100000100001100100110001",
3025 => "0101000100000100100100011",
3026 => "0100000001010010011110001",
3027 => "0101100001000110011100011",
3028 => "0011001011001100011010001",
3029 => "0100101011000110011000010",
3030 => "0111001100001000101110001",
3031 => "0111001100000100101100010",
3032 => "0011001100001000101110001",
3033 => "0100001100000100101100010",
3034 => "0100000000011001001010001",
3035 => "0110000000001001001000011",
3036 => "0001001100010100010110001",
3037 => "0011101100001010010100010",
3038 => "0001010100101100001110001",
3039 => "0001010101101100000100011",
3040 => "0000000100000101010010001",
3041 => "0000100100000011010000010",
3042 => "0000000010110000010010001",
3043 => "0100000010010000010000011",
3044 => "0011101000010100010010001",
3045 => "0011101010010100001000010",
3046 => "0011000111010000101010001",
3047 => "0011000111001000010100010",
3048 => "0101001100001000010100010",
3049 => "0111000000001100111010001",
3050 => "1000100000000110011100010",
3051 => "0111000111000110011100010",
3052 => "0010001011001010100010001",
3053 => "0010001111001010010000010",
3054 => "0001000000101000100110001",
3055 => "0001000011101000001100011",
3056 => "0011000111011000100010001",
3057 => "0011000111001100010000010",
3058 => "0110001011001100010000010",
3059 => "0100110001001100011010001",
3060 => "0100110100001100001100010",
3061 => "0011101010010100010010001",
3062 => "0011101100010100001000010",
3063 => "0011000101011000100110001",
3064 => "0101000101001000100100011",
3065 => "0010101011001100100010001",
3066 => "0100001011000110100000010",
3067 => "1001000100001001000110001",
3068 => "1001000100000101000100010",
3069 => "0000000000001100011010001",
3070 => "0001100000000110011000010",
3071 => "1001000100001001000110001",
3072 => "1001000100000101000100010",
3073 => "0001000100001001000110001",
3074 => "0010000100000101000100010",
3075 => "0010110010100110001110001",
3076 => "0010110011100110000100011",
3077 => "0101100000000101001010001",
3078 => "0101101001000100100100010",
3079 => "0111100100000101001010001",
3080 => "0111101101000100100100010",
3081 => "0011100100000101001010001",
3082 => "0011101101000100100100010",
3083 => "0011101011010100100010001",
3084 => "0110001011001010010000010",
3085 => "0011101111001010010000010",
3086 => "0101000110001000100110001",
3087 => "0110000110000100100100010",
3088 => "0101000000001100100110001",
3089 => "0110000000000100100100011",
3090 => "0001001001100000100010001",
3091 => "0001001001010000010000010",
3092 => "0101001101010000010000010",
3093 => "0111001111001100100110001",
3094 => "0111010010001100001100011",
3095 => "0100000111001100100110001",
3096 => "0101000111000100100100011",
3097 => "0111001111001100100110001",
3098 => "0111010010001100001100011",
3099 => "0001101100011000011010001",
3100 => "0001101110011000001000011",
3101 => "0111001100010010011010001",
3102 => "0111001110010010001000011",
3103 => "0000101100010010011010001",
3104 => "0000101110010010001000011",
3105 => "0001100111100100001110001",
3106 => "0001101000100100000100011",
3107 => "0000100111101100011010001",
3108 => "0000101001101100001000011",
3109 => "1001000100001100011010001",
3110 => "1001000111001100001100010",
3111 => "0000000100001100011010001",
3112 => "0000000111001100001100010",
3113 => "0010101011100000011010001",
3114 => "0010101110100000001100010",
3115 => "0011010000010010010010001",
3116 => "0011010010010010001000010",
3117 => "0111001111001100100110001",
3118 => "0111010010001100001100011",
3119 => "0010001111001100100110001",
3120 => "0010010010001100001100011",
3121 => "0111100001001101011110001",
3122 => "1000100001000101011100011",
3123 => "0000010101110000001110001",
3124 => "0100010101010000001100011",
3125 => "0000010100110000010010001",
3126 => "0100010100010000010000011",
3127 => "0001100001001101011110001",
3128 => "0010100001000101011100011",
3129 => "0001110001100100001110001",
3130 => "0001110010100100000100011",
3131 => "0000010000100100001110001",
3132 => "0000010001100100000100011",
3133 => "0000110000101100010010001",
3134 => "0110010000010110001000010",
3135 => "0000110010010110001000010",
3136 => "0000010000010010011010001",
3137 => "0000010010010010001000011",
3138 => "0001001010101010001110001",
3139 => "0100101010001110001100011",
3140 => "0001010010011000011010001",
3141 => "0001010010001100001100010",
3142 => "0100010101001100001100010",
3143 => "0000000101110000010010001",
3144 => "0000000111110000001000010",
3145 => "0101000010001000111110001",
3146 => "0101000111001000010100011",
3147 => "0101000111001100110010001",
3148 => "0101001101001100011000010",
3149 => "0011000110001100100110001",
3150 => "0100000110000100100100011",
3151 => "0101100000001100100110001",
3152 => "0110100000000100100100011",
3153 => "0100100111001100100110001",
3154 => "0101100111000100100100011",
3155 => "0001000001101000001110001",
3156 => "0001000010101000000100011",
3157 => "0000110010011000011010001",
3158 => "0000110010001100001100010",
3159 => "0011110101001100001100010",
3160 => "0110100010001000110110001",
3161 => "0110100010000100110100010",
3162 => "0011000111011000010010001",
3163 => "0110000111001100010000010",
3164 => "0101000001001000110110001",
3165 => "0101000001000100110100010",
3166 => "0011000000000111001010001",
3167 => "0011100000000011001000011",
3168 => "0111000011010100010110001",
3169 => "0111000011001010010100010",
3170 => "0011001111011000100010001",
3171 => "0101001111001000100000011",
3172 => "0100101010001100100110001",
3173 => "0101101010000100100100011",
3174 => "0100000011001000100110001",
3175 => "0101000011000100100100010",
3176 => "1000100000001100111010001",
3177 => "1010000000000110011100010",
3178 => "1000100111000110011100010",
3179 => "0000100000001100111010001",
3180 => "0000100000000110011100010",
3181 => "0010000111000110011100010",
3182 => "0111000000001101000010001",
3183 => "1000100000000110100000010",
3184 => "0111001000000110100000010",
3185 => "0011100100001000101010001",
3186 => "0100100100000100101000010",
3187 => "0001110001100100011010001",
3188 => "0110010001010010001100010",
3189 => "0001110100010010001100010",
3190 => "0000110100101100010010001",
3191 => "0110010100010110010000010",
3192 => "0111000011010100010110001",
3193 => "0111000011001010010100010",
3194 => "0000000011010100010110001",
3195 => "0010100011001010010100010",
3196 => "0110000110011001000010001",
3197 => "1000000110001001000000011",
3198 => "0000000110011001000010001",
3199 => "0010000110001001000000011",
3200 => "0101001001001010111110001",
3201 => "0101001110001010010100011",
3202 => "0000110010101010001010001",
3203 => "0000110011101010000100010",
3204 => "0111100000010010011010001",
3205 => "0111100010010010001000011",
3206 => "0011000001011000010010001",
3207 => "0110000001001100010000010",
3208 => "0011000000011000110010001",
3209 => "0110000000001100011000010",
3210 => "0011000110001100011000010",
3211 => "0100001010010000110010001",
3212 => "0100001010001000011000010",
3213 => "0110010000001000011000010",
3214 => "0111010000010100100010001",
3215 => "1001110000001010010000010",
3216 => "0111010100001010010000010",
3217 => "0000010000010100100010001",
3218 => "0000010000001010010000010",
3219 => "0010110100001010010000010",
3220 => "0101001100011000010110001",
3221 => "0111001100001000010100011",
3222 => "0011010000010100100010001",
3223 => "0011010000001010010000010",
3224 => "0101110100001010010000010",
3225 => "0011100110011000011010001",
3226 => "0110100110001100001100010",
3227 => "0011101001001100001100010",
3228 => "0100100110001001001010001",
3229 => "0100100110000100100100010",
3230 => "0101101111000100100100010",
3231 => "0101001001001100111010001",
3232 => "0110101001000110011100010",
3233 => "0101010000000110011100010",
3234 => "0100001001001100111010001",
3235 => "0100001001000110011100010",
3236 => "0101110000000110011100010",
3237 => "0011100100010110110010001",
3238 => "0011101010010110011000010",
3239 => "0010001000001101000010001",
3240 => "0010001000000110100000010",
3241 => "0011110000000110100000010",
3242 => "1000100011001001010110001",
3243 => "1000101010001000011100011",
3244 => "0001100011001001010110001",
3245 => "0001101010001000011100011",
3246 => "0101000001010001001010001",
3247 => "0111000001001000100100010",
3248 => "0101001010001000100100010",
3249 => "0001000101100000100010001",
3250 => "0001000101010000010000010",
3251 => "0101001001010000010000010",
3252 => "0001100110100100110010001",
3253 => "0001101010100100010000011",
3254 => "0010001010100000110010001",
3255 => "0010001110100000010000011",
3256 => "0111100100010001010010001",
3257 => "1001100100001000101000010",
3258 => "0111101110001000101000010",
3259 => "0011100010010010011010001",
3260 => "0101000010000110011000011",
3261 => "0111100100010001010010001",
3262 => "1001100100001000101000010",
3263 => "0111101110001000101000010",
3264 => "0000100100010001010010001",
3265 => "0000100100001000101000010",
3266 => "0010101110001000101000010",
3267 => "0101101000010000111010001",
3268 => "0111101000001000011100010",
3269 => "0101101111001000011100010",
3270 => "0010101000010000111010001",
3271 => "0010101000001000011100010",
3272 => "0100101111001000011100010",
3273 => "0101001101001010100010001",
3274 => "0101010001001010010000010",
3275 => "0010001101001110100110001",
3276 => "0010010000001110001100011",
3277 => "0000001101110000101010001",
3278 => "0000010010110000010100010",
3279 => "0010000010010000101110001",
3280 => "0100000010001000101100010",
3281 => "0101000010010001000010001",
3282 => "0111000010001000100000010",
3283 => "0101001010001000100000010",
3284 => "0000000010110000011010001",
3285 => "0000000010011000001100010",
3286 => "0110000101011000001100010",
3287 => "0011000000011000100110001",
3288 => "0011000011011000001100011",
3289 => "0000100010011000110010001",
3290 => "0000100010001100011000010",
3291 => "0011101000001100011000010",
3292 => "1001000101001100100110001",
3293 => "1001001000001100001100011",
3294 => "0010000011010000101010001",
3295 => "0010000011001000010100010",
3296 => "0100001000001000010100010",
3297 => "0011010101100100001110001",
3298 => "0011010110100100000100011",
3299 => "0000101010100100001010001",
3300 => "0000101011100100000100010",
3301 => "0000101010101100001110001",
3302 => "0000101011101100000100011",
3303 => "0001001000011000100110001",
3304 => "0001001011011000001100011",
3305 => "0110001000011000011010001",
3306 => "1001001000001100001100010",
3307 => "0110001011001100001100010",
3308 => "0000001000011000011010001",
3309 => "0000001000001100001100010",
3310 => "0011001011001100001100010",
3311 => "0101001111001100100110001",
3312 => "0110001111000100100100011",
3313 => "0011101101010010011010001",
3314 => "0011101111010010001000011",
3315 => "0100101000001110110010001",
3316 => "0100101110001110011000010",
3317 => "0010001101010010011010001",
3318 => "0011101101000110011000011",
3319 => "0011001111100100010010001",
3320 => "0110001111001100010000011",
3321 => "0010100100001001000010001",
3322 => "0011100100000101000000010",
3323 => "0101001111001100100110001",
3324 => "0110001111000100100100011",
3325 => "0100001111001100100110001",
3326 => "0101001111000100100100011",
3327 => "0100101011011000101010001",
3328 => "0111101011001100010100010",
3329 => "0100110000001100010100010",
3330 => "0001100110011100011010001",
3331 => "0001101000011100001000011",
3332 => "0010000010100010100010001",
3333 => "0010000110100010010000010",
3334 => "0011000010011001010110001",
3335 => "0011001001011000011100011",
3336 => "0100000001010010100110001",
3337 => "0100000100010010001100011",
3338 => "0000000111110000001110001",
3339 => "0110000111011000001100010",
3340 => "0101100110010010101010001",
3341 => "0101101011010010010100010",
3342 => "0001001011100100001110001",
3343 => "0001001100100100000100011",
3344 => "0100010000010010010010001",
3345 => "0100010010010010001000010",
3346 => "0000000000010010011010001",
3347 => "0000000010010010001000011",
3348 => "0000001011110000011010001",
3349 => "0000001101110000001000011",
3350 => "0001001001101000011010001",
3351 => "0001001100101000001100010",
3352 => "0010000101100000110010001",
3353 => "0110000101010000011000010",
3354 => "0010001011010000011000010",
3355 => "0101000010001000111110001",
3356 => "0101000111001000010100011",
3357 => "0011100011010100010010001",
3358 => "0011100101010100001000010",
3359 => "0100101111001100100010001",
3360 => "0100110011001100010000010",
3361 => "1000100000001110101010001",
3362 => "1000100101001110010100010",
3363 => "0000000000001110101010001",
3364 => "0000000101001110010100010",
3365 => "1000000001001100110010001",
3366 => "1001100001000110011000010",
3367 => "1000000111000110011000010",
3368 => "0000100000100110100010001",
3369 => "0000100100100110010000010",
3370 => "0110000010010010010010001",
3371 => "0110000100010010001000010",
3372 => "0001100010010010010010001",
3373 => "0001100100010010001000010",
3374 => "0110000010010100011010001",
3375 => "0110000100010100001000011",
3376 => "0001100100100100001010001",
3377 => "0110000100010010001000010",
3378 => "0110000001001000100110001",
3379 => "0110000001000100100100010",
3380 => "0100000001001000100110001",
3381 => "0101000001000100100100010",
3382 => "0101000101010000101010001",
3383 => "0111000101001000010100010",
3384 => "0101001010001000010100010",
3385 => "0011000100011000110110001",
3386 => "0101000100001000110100011",
3387 => "0110100101001100011010001",
3388 => "0110100101000110011000010",
3389 => "0000100101011000001110001",
3390 => "0011100101001100001100010",
3391 => "0011100101010100011010001",
3392 => "0011100111010100001000011",
3393 => "0001000000101010010110001",
3394 => "0100100000001110010100011",
3395 => "0000001000010010100110001",
3396 => "0000001011010010001100011",
3397 => "0100100110001100100110001",
3398 => "0101100110000100100100011",
3399 => "0000000011001100011110001",
3400 => "0001100011000110011100010",
3401 => "0100110010011000011010001",
3402 => "0111110010001100001100010",
3403 => "0100110101001100001100010",
3404 => "0001001000101000011010001",
3405 => "0001001000010100001100010",
3406 => "0110001011010100001100010",
3407 => "0110100010010100010010001",
3408 => "0110100100010100001000010",
3409 => "0010000101001011001010001",
3410 => "0010001011001010011000011",
3411 => "1010000100001000100110001",
3412 => "1010000100000100100100010",
3413 => "0100000110010000111010001",
3414 => "0100001101010000011100010",
3415 => "0000000001110000011010001",
3416 => "0110000001011000001100010",
3417 => "0000000100011000001100010",
3418 => "0000000100001000100110001",
3419 => "0001000100000100100100010",
3420 => "0001100110100100001110001",
3421 => "0001100111100100000100011",
3422 => "0001110001100000011010001",
3423 => "0001110011100000001000011",
3424 => "0110100110001100100110001",
3425 => "0110101001001100001100011",
3426 => "0010100110011100011010001",
3427 => "0010100110001110001100010",
3428 => "0110001001001110001100010",
3429 => "0110100101010000101010001",
3430 => "1000100101001000010100010",
3431 => "0110101010001000010100010",
3432 => "0001000010101000001110001",
3433 => "0001000011101000000100011",
3434 => "0100100010010010011010001",
3435 => "0110000010000110011000011",
3436 => "0100000110001100100110001",
3437 => "0101000110000100100100011",
3438 => "0110000011001000101110001",
3439 => "0110000011000100101100010",
3440 => "0100000011001000101110001",
3441 => "0101000011000100101100010",
3442 => "0100000011010000101010001",
3443 => "0110000011001000010100010",
3444 => "0100001000001000010100010",
3445 => "0101100001000101001010001",
3446 => "0110000001000011001000010",
3447 => "0100100010010010011010001",
3448 => "0110000010000110011000011",
3449 => "0000000010100110001110001",
3450 => "0000000011100110000100011",
3451 => "0100101110010010011010001",
3452 => "0100110000010010001000011",
3453 => "0000101000100100010110001",
3454 => "0011101000001100010100011",
3455 => "0110000000001100100110001",
3456 => "0111000000000100100100011",
3457 => "0011000000001100100110001",
3458 => "0100000000000100100100011",
3459 => "0110100110001000111110001",
3460 => "0110101011001000010100011",
3461 => "0000100101100100001110001",
3462 => "0000100110100100000100011",
3463 => "0100100111011100011010001",
3464 => "0100101001011100001000011",
3465 => "0001010000100100001110001",
3466 => "0001010001100100000100011",
3467 => "0111110001010010011010001",
3468 => "0111110011010010001000011",
3469 => "0000001000011000011010001",
3470 => "0000001000001100001100010",
3471 => "0011001011001100001100010",
3472 => "0100101101001110100010001",
3473 => "0100110001001110010000010",
3474 => "0001010001101000001110001",
3475 => "0001010010101000000100011",
3476 => "0111110001010010011010001",
3477 => "0111110011010010001000011",
3478 => "0010000000011110010010001",
3479 => "0010000010011110001000010",
3480 => "1000100010001100011010001",
3481 => "1000100101001100001100010",
3482 => "0000000011001100100110001",
3483 => "0000000110001100001100011",
3484 => "0111110001010010011010001",
3485 => "0111110011010010001000011",
3486 => "0000010001010010011010001",
3487 => "0000010011010010001000011",
3488 => "0100110010011000011010001",
3489 => "0111110010001100001100010",
3490 => "0100110101001100001100010",
3491 => "0001101111001100100110001",
3492 => "0001110010001100001100011",
3493 => "1000001101010000101010001",
3494 => "1010001101001000010100010",
3495 => "1000010010001000010100010",
3496 => "0000001110110000010010001",
3497 => "0100001110010000010000011",
3498 => "0110110010001100011010001",
3499 => "0110110010000110011000010",
3500 => "0000001101010000101010001",
3501 => "0000001101001000010100010",
3502 => "0010010010001000010100010",
3503 => "0000001110110000011010001",
3504 => "0000010001110000001100010",
3505 => "0010100010011000100010001",
3506 => "0010100010001100010000010",
3507 => "0101100110001100010000010",
3508 => "0100001001010010011010001",
3509 => "0101101001000110011000011",
3510 => "0010000011100000010010001",
3511 => "0010000101100000001000010",
3512 => "0101000010001000101010001",
3513 => "0101000111001000010100010",
3514 => "0100000100001010100010001",
3515 => "0100001000001010010000010",
3516 => "0101100101010010110010001",
3517 => "0101101001010010010000011",
3518 => "0010000101010010110010001",
3519 => "0010001001010010010000011",
3520 => "0111000110001100100110001",
3521 => "0111001001001100001100011",
3522 => "0001000100101000110010001",
3523 => "0001001000101000010000011",
3524 => "0010000100100011000010001",
3525 => "0010001100100010100000010",
3526 => "0100000111001110011010001",
3527 => "0100001010001110001100010",
3528 => "0000101001101110001010001",
3529 => "0000101010101110000100010",
3530 => "0011100000001100100110001",
3531 => "0100100000000100100100011",
3532 => "0110100011001000100110001",
3533 => "0110100011000100100100010",
3534 => "0100000001001100110110001",
3535 => "0101000001000100110100011",
3536 => "0010010110100100001010001",
3537 => "0010010111100100000100010",
3538 => "0001101010010010011010001",
3539 => "0011001010000110011000011",
3540 => "0111000000000101100010001",
3541 => "0111000000000011100000010",
3542 => "0100000000000101100010001",
3543 => "0100100000000011100000010",
3544 => "0001100010100100101010001",
3545 => "0100100010001100101000011",
3546 => "0010001101011110011010001",
3547 => "0100101101001010011000011",
3548 => "0001110101100100001110001",
3549 => "0100110101001100001100011",
3550 => "0100100001001000101110001",
3551 => "0101100001000100101100010",
3552 => "0100100111010100010010001",
3553 => "0100100111001010010000010",
3554 => "0011100000010101001010001",
3555 => "0110000000001011001000010",
3556 => "0110000001001101000010001",
3557 => "0111000001000101000000011",
3558 => "0011000001001101000010001",
3559 => "0100000001000101000000011",
3560 => "1001000010001100011010001",
3561 => "1001000101001100001100010",
3562 => "0001100101100100001010001",
3563 => "0001100110100100000100010",
3564 => "1001000010001100011010001",
3565 => "1001000101001100001100010",
3566 => "0000000010001100011010001",
3567 => "0000000101001100001100010",
3568 => "0110101011010110011010001",
3569 => "0110101101010110001000011",
3570 => "0010100111010100010010001",
3571 => "0101000111001010010000010",
3572 => "0101101001010100011110001",
3573 => "0101101001001010011100010",
3574 => "0001101001010100011110001",
3575 => "0100001001001010011100010",
3576 => "1000000100001100011010001",
3577 => "1000000100000110011000010",
3578 => "0010100110010100100010001",
3579 => "0010100110001010010000010",
3580 => "0101001010001010010000010",
3581 => "0011110101100000001110001",
3582 => "0011110101010000001100010",
3583 => "0000110101100000001110001",
3584 => "0100110101010000001100010",
3585 => "0001000101101100111010001",
3586 => "0110100101010110011100010",
3587 => "0001001100010110011100010",
3588 => "0001101010010000101010001",
3589 => "0001101010001000010100010",
3590 => "0011101111001000010100010",
3591 => "1000100000001100110010001",
3592 => "1010000000000110011000010",
3593 => "1000100110000110011000010",
3594 => "0010100010001101001010001",
3595 => "0011100010000101001000011",
3596 => "0110100000001100100110001",
3597 => "0111100000000100100100011",
3598 => "0000001100001110100110001",
3599 => "0000001111001110001100011",
3600 => "0111101101010000101010001",
3601 => "1001101101001000010100010",
3602 => "0111110010001000010100010",
3603 => "0000100000001100110010001",
3604 => "0000100000000110011000010",
3605 => "0010000110000110011000010",
3606 => "0110000001000110110010001",
3607 => "0110000111000110011000010",
3608 => "0000101101010000101010001",
3609 => "0000101101001000010100010",
3610 => "0010110010001000010100010",
3611 => "0001110101100110001010001",
3612 => "0001110110100110000100010",
3613 => "0011000011001000110110001",
3614 => "0100000011000100110100010",
3615 => "0010101010100100001110001",
3616 => "0010101011100100000100011",
3617 => "0100100011001010110010001",
3618 => "0100100111001010010000011",
3619 => "0101100010001000111110001",
3620 => "0101100111001000010100011",
3621 => "0010000001100000010010001",
3622 => "0010000011100000001000010",
3623 => "0011000000100100001110001",
3624 => "0011000001100100000100011",
3625 => "0010100001010100100010001",
3626 => "0010100001001010010000010",
3627 => "0101000101001010010000010",
3628 => "0101110010011000011010001",
3629 => "1000110010001100001100010",
3630 => "0101110101001100001100010",
3631 => "0010101111011000001110001",
3632 => "0101101111001100001100010",
3633 => "0000101010101100010010001",
3634 => "0000101010010110010000010",
3635 => "0011101001010010011010001",
3636 => "0101001001000110011000011",
3637 => "0011001011011000010110001",
3638 => "0101001011001000010100011",
3639 => "0011000111010100011110001",
3640 => "0101100111001010011100010",
3641 => "0101100010010000101010001",
3642 => "0101100010001000101000010",
3643 => "0010100010010000101010001",
3644 => "0100100010001000101000010",
3645 => "0011000100100100011010001",
3646 => "0111100100010010001100010",
3647 => "0011000111010010001100010",
3648 => "0000000101010100100110001",
3649 => "0000001000010100001100011",
3650 => "0001000111101010011010001",
3651 => "0001001001101010001000011",
3652 => "0000000100101101000010001",
3653 => "0000000100010110100000010",
3654 => "0101101100010110100000010",
3655 => "0100100000001101011010001",
3656 => "0100101011001100101100010",
3657 => "0100100001000110110010001",
3658 => "0100100111000110011000010",
3659 => "0110000000011001001010001",
3660 => "1001000000001100100100010",
3661 => "0110001001001100100100010",
3662 => "0000000000011001001010001",
3663 => "0000000000001100100100010",
3664 => "0011001001001100100100010",
3665 => "0000100001101100010010001",
3666 => "0110000001010110001000010",
3667 => "0000100011010110001000010",
3668 => "0001100000100100010010001",
3669 => "0001100010100100001000010",
3670 => "0001000101101100011010001",
3671 => "0001000111101100001000011",
3672 => "0010100000001100100110001",
3673 => "0010100011001100001100011",
3674 => "0101001110001100100110001",
3675 => "0110001110000100100100011",
3676 => "0100001110001100100110001",
3677 => "0101001110000100100100011",
3678 => "0010110010100100001110001",
3679 => "0010110011100100000100011",
3680 => "0011000000001100110110001",
3681 => "0100100000000110110100010",
3682 => "0011100100011000010010001",
3683 => "0011100100001100010000010",
3684 => "0010100010011000011010001",
3685 => "0100100010001000011000011",
3686 => "0010000001100100001110001",
3687 => "0010000010100100000100011",
3688 => "0000001000001100110010001",
3689 => "0000001100001100010000011",
3690 => "0100101111001100100110001",
3691 => "0101101111000100100100011",
3692 => "0100101010001100110110001",
3693 => "0101101010000100110100011",
3694 => "0011010001100100001010001",
3695 => "0011010010100100000100010",
3696 => "0100100100001100100110001",
3697 => "0101100100000100100100011",
3698 => "0101000000001100100110001",
3699 => "0110000000000100100100011",
3700 => "0010100110010100100010001",
3701 => "0010100110001010010000010",
3702 => "0101001010001010010000010",
3703 => "0111001001001010100010001",
3704 => "0111001101001010010000010",
3705 => "0010101001001010100010001",
3706 => "0010101101001010010000010",
3707 => "0111001011010010011010001",
3708 => "0111001101010010001000011",
3709 => "0000000010101110111110001",
3710 => "0000000111101110010100011",
3711 => "1000000000010000110010001",
3712 => "1000000110010000011000010",
3713 => "0010001111001100100110001",
3714 => "0010010010001100001100011",
3715 => "0100010010010010010010001",
3716 => "0100010100010010001000010",
3717 => "0000010001100100001110001",
3718 => "0000010010100100000100011",
3719 => "0110101011010110011010001",
3720 => "0110101101010110001000011",
3721 => "0000001011010110011010001",
3722 => "0000001101010110001000011",
3723 => "0000001001110000011010001",
3724 => "0110001001011000001100010",
3725 => "0000001100011000001100010",
3726 => "0011010000010000100010001",
3727 => "0011010100010000010000010",
3728 => "0101010000011100011010001",
3729 => "0101010010011100001000011",
3730 => "0000100001101010001110001",
3731 => "0000100010101010000100011",
3732 => "0000000010110000001110001",
3733 => "0000000010011000001100010",
3734 => "0001001111010000010110001",
3735 => "0011001111001000010100010",
3736 => "0001001011101010001110001",
3737 => "0100101011001110001100011",
3738 => "0000110010011000011010001",
3739 => "0000110010001100001100010",
3740 => "0011110101001100001100010",
3741 => "0101001110001000101010001",
3742 => "0101010011001000010100010",
3743 => "0011100111001000101010001",
3744 => "0011101100001000010100010",
3745 => "0100101000001100110010001",
3746 => "0100101100001100010000011",
3747 => "0011100001010010011010001",
3748 => "0101000001000110011000011",
3749 => "0001101110100110001010001",
3750 => "0001101111100110000100010",
3751 => "0011100111010100101010001",
3752 => "0011100111001010010100010",
3753 => "0110001100001010010100010",
3754 => "0001101100100100110010001",
3755 => "0001101100010010110000010",
3756 => "0100000000001100110010001",
3757 => "0101000000000100110000011",
3758 => "0001100000100010100110001",
3759 => "0001100011100010001100011",
3760 => "0011000000011000101110001",
3761 => "0101000000001000101100011",
3762 => "0000100000001100110110001",
3763 => "0010000000000110110100010",
3764 => "0010101000100000011010001",
3765 => "0010101011100000001100010",
3766 => "0100001000001010110010001",
3767 => "0100001110001010011000010",
3768 => "0001110101100100001110001",
3769 => "0100110101001100001100011",
3770 => "0000000000001100011010001",
3771 => "0001100000000110011000010",
3772 => "0001000000101000001110001",
3773 => "0001000001101000000100011",
3774 => "0010000110011110101010001",
3775 => "0100100110001010101000011",
3776 => "0100100110001100100110001",
3777 => "0101100110000100100100011",
3778 => "0100100000001100100110001",
3779 => "0101100000000100100100011",
3780 => "0111000000001100100110001",
3781 => "1000000000000100100100011",
3782 => "0011110000010010011010001",
3783 => "0011110010010010001000011",
3784 => "0111000000001100100110001",
3785 => "1000000000000100100100011",
3786 => "0010000000001100100110001",
3787 => "0011000000000100100100011",
3788 => "1000100001001101000010001",
3789 => "1001100001000101000000011",
3790 => "0000100001001101000010001",
3791 => "0001100001000101000000011",
3792 => "0111001101001100100110001",
3793 => "0111010000001100001100011",
3794 => "0000000000001100100110001",
3795 => "0000000011001100001100011",
3796 => "0100100101001100011010001",
3797 => "0100100101000110011000010",
3798 => "0001101010010010011010001",
3799 => "0011001010000110011000011",
3800 => "0111000111000111000010001",
3801 => "0111001111000110100000010",
3802 => "0010001010011100110010001",
3803 => "0010001010001110011000010",
3804 => "0101110000001110011000010",
3805 => "0011100110011000011010001",
3806 => "0011101000011000001000011",
3807 => "0011100010001001010010001",
3808 => "0100100010000101010000010",
3809 => "0111001101001100100110001",
3810 => "0111010000001100001100011",
3811 => "0101000110001000100110001",
3812 => "0110000110000100100100010",
3813 => "0111001101001100100110001",
3814 => "0111010000001100001100011",
3815 => "0010110100011100010010001",
3816 => "0010110110011100001000010",
3817 => "0010000100100000110010001",
3818 => "0010001010100000011000010",
3819 => "0100100110001100100110001",
3820 => "0101100110000100100100011",
3821 => "0001100000101010010010001",
3822 => "0001100010101010001000010",
3823 => "0010001101001100100110001",
3824 => "0010010000001100001100011",
3825 => "1000010000001010100010001",
3826 => "1000010100001010010000010",
3827 => "0010000000100001000010001",
3828 => "0010000000010000100000010",
3829 => "0110001000010000100000010",
3830 => "0011000110011100011010001",
3831 => "0110100110001110001100010",
3832 => "0011001001001110001100010",
3833 => "0101000101001000111110001",
3834 => "0101001010001000010100011",
3835 => "0100101111011000100010001",
3836 => "0111101111001100010000010",
3837 => "0100110011001100010000010",
3838 => "0011000111011000010010001",
3839 => "0110000111001100010000010",
3840 => "0010100110011100011010001",
3841 => "0110000110001110001100010",
3842 => "0010101001001110001100010",
3843 => "0001100110100100101010001",
3844 => "0001100110010010010100010",
3845 => "0110001011010010010100010",
3846 => "0011000000100101010110001",
3847 => "0110000000001101010100011",
3848 => "0000000000110001010110001",
3849 => "0100000000010001010100011",
3850 => "0011010010100100001110001",
3851 => "0011010011100100000100011",
3852 => "0000001111010010011010001",
3853 => "0000010001010010001000011",
3854 => "0010000011100110001010001",
3855 => "0010000100100110000100010",
3856 => "0000000011110000001010001",
3857 => "0000000100110000000100010",
3858 => "0111101110010010010010001",
3859 => "0111110000010010001000010",
3860 => "0000001110010010010010001",
3861 => "0000010000010010001000010",
3862 => "0011001111100100001010001",
3863 => "0011010000100100000100010",
3864 => "0001110001100100001110001",
3865 => "0001110010100100000100011",
3866 => "0110000000000111011110001",
3867 => "0110100000000011011100011",
3868 => "0011000000010000011010001",
3869 => "0011000011010000001100010",
3870 => "0011010000100100001110001",
3871 => "0011010001100100000100011",
3872 => "0100100000000111011110001",
3873 => "0101000000000011011100011",
3874 => "0101000111001000101010001",
3875 => "0101001100001000010100010",
3876 => "0011101000010100110010001",
3877 => "0011101100010100010000011",
3878 => "0111001001001100111010001",
3879 => "1000101001000110011100010",
3880 => "0111010000000110011100010",
3881 => "0001000000010100100110001",
3882 => "0001000011010100001100011",
3883 => "0101100001001010110010001",
3884 => "0101100111001010011000010",
3885 => "0000100100011000101010001",
3886 => "0000100100001100010100010",
3887 => "0011101001001100010100010",
3888 => "0111100001010010010010001",
3889 => "0111100011010010001000010",
3890 => "0000100010010000101010001",
3891 => "0000100010001000010100010",
3892 => "0010100111001000010100010",
3893 => "0101000001001010110010001",
3894 => "0101000101001010010000011",
3895 => "0010000000011101100010001",
3896 => "0101100000001111100000010",
3897 => "0011110001010100010010001",
3898 => "0011110011010100001000010",
3899 => "0101001110001000101010001",
3900 => "0101010011001000010100010",
3901 => "0110101111001100100110001",
3902 => "0111101111000100100100011",
3903 => "0001110101100100001110001",
3904 => "0001110110100100000100011",
3905 => "0110101111001100100110001",
3906 => "0111101111000100100100011",
3907 => "0010101111001100100110001",
3908 => "0011101111000100100100011",
3909 => "0101000110001001001010001",
3910 => "0110000110000100100100010",
3911 => "0101001111000100100100010",
3912 => "0011100011001100101110001",
3913 => "0100100011000100101100011",
3914 => "0111100001010010010010001",
3915 => "0111100011010010001000010",
3916 => "0010100100011100100010001",
3917 => "0010101000011100010000010",
3918 => "0100000001011110100110001",
3919 => "0100000100011110001100011",
3920 => "0011100010010000101010001",
3921 => "0011100010001000010100010",
3922 => "0101100111001000010100010",
3923 => "0110000010001100110010001",
3924 => "0110000010000110110000010",
3925 => "0011000010001100110010001",
3926 => "0100100010000110110000010",
3927 => "0011100111011000010010001",
3928 => "0011100111001100010000010",
3929 => "0011000011011000101010001",
3930 => "0101000011001000101000011",
3931 => "0010100110100000011010001",
3932 => "0110100110010000001100010",
3933 => "0010101001010000001100010",
3934 => "0001100001100100100110001",
3935 => "0100100001001100100100011",
3936 => "0001101000100100010110001",
3937 => "0100101000001100010100011",
3938 => "0000000000110001011010001",
3939 => "0000000000011000101100010",
3940 => "0110001011011000101100010",
3941 => "0111010000010010011010001",
3942 => "0111010010010010001000011",
3943 => "0000010000110000100010001",
3944 => "0000010100110000010000010",
3945 => "0000110011101100010010001",
3946 => "0110010011010110001000010",
3947 => "0000110101010110001000010",
3948 => "0000110000010010011010001",
3949 => "0000110010010010001000011",
3950 => "0011101000010100010010001",
3951 => "0011101000001010010000010",
3952 => "0100101111001100100110001",
3953 => "0101101111000100100100011",
3954 => "0101010010011000011010001",
3955 => "1000010010001100001100010",
3956 => "0101010101001100001100010",
3957 => "0001010010011000011010001",
3958 => "0001010010001100001100010",
3959 => "0100010101001100001100010",
3960 => "0100000011100000100110001",
3961 => "0100000110100000001100011",
3962 => "0000000101010100011010001",
3963 => "0000000111010100001000011",
3964 => "0010100101100100001110001",
3965 => "0010100110100100000100011",
3966 => "0001000110010010011010001",
3967 => "0001001001010010001100010",
3968 => "0111000010010100100110001",
3969 => "0111000101010100001100011",
3970 => "0001100110100100001110001",
3971 => "0001100111100100000100011",
3972 => "0100100010011110011010001",
3973 => "0100100100011110001000011",
3974 => "0010001000011110011010001",
3975 => "0010001010011110001000011",
3976 => "0000000101110000010010001",
3977 => "0110000101011000001000010",
3978 => "0000000111011000001000010",
3979 => "0011101000001100110010001",
3980 => "0100101000000100110000011",
3981 => "0101100000001100100110001",
3982 => "0110100000000100100100011",
3983 => "0000001100001100110010001",
3984 => "0000001100000110011000010",
3985 => "0001110010000110011000010",
3986 => "0111001100010100011010001",
3987 => "0111001110010100001000011",
3988 => "0001000111100100100110001",
3989 => "0001001010100100001100011",
3990 => "0101101110010100100110001",
3991 => "0101110001010100001100011",
3992 => "0011100110010100100010001",
3993 => "0011100110001010010000010",
3994 => "0110001010001010010000010",
3995 => "0011000110011100011010001",
3996 => "0110100110001110001100010",
3997 => "0011001001001110001100010",
3998 => "0010001101010010011110001",
3999 => "0011101101000110011100011",
4000 => "0111001010001100110010001",
4001 => "1000101010000110011000010",
4002 => "0111010000000110011000010",
4003 => "0010001010001100110010001",
4004 => "0010001010000110011000010",
4005 => "0011110000000110011000010",
4006 => "0110101001010000011010001",
4007 => "0110101001001000011000010",
4008 => "0100000011001000111010001",
4009 => "0101000011000100111000010",
4010 => "1000100000000111001010001",
4011 => "1001000000000011001000011",
4012 => "0010001100100000110010001",
4013 => "0110001100010000110000010",
4014 => "0111100000001100111010001",
4015 => "1000100000000100111000011",
4016 => "0001100000001100111010001",
4017 => "0010100000000100111000011",
4018 => "0110000010011001010010001",
4019 => "1000000010001001010000011",
4020 => "0000000010011001010010001",
4021 => "0010000010001001010000011",
4022 => "1000000000001101000110001",
4023 => "1001000000000101000100011",
4024 => "0001000000001101000110001",
4025 => "0010000000000101000100011",
4026 => "0111100110010010011010001",
4027 => "0111101000010010001000011",
4028 => "0000000110010010011010001",
4029 => "0000001000010010001000011",
4030 => "1001000001001100110110001",
4031 => "1010000001000100110100011",
4032 => "0000000001001100110110001",
4033 => "0001000001000100110100011",
4034 => "1000000000001000100110001",
4035 => "1000000000000100100100010",
4036 => "0010101010011000011110001",
4037 => "0100101010001000011100011",
4038 => "0110001001011000011010001",
4039 => "0110001011011000001000011",
4040 => "0000001001011000011010001",
4041 => "0000001011011000001000011",
4042 => "0010100111011100100110001",
4043 => "0010101010011100001100011",
4044 => "0000001111101000001110001",
4045 => "0000010000101000000100011",
4046 => "0100001010010000101010001",
4047 => "0110001010001000010100010",
4048 => "0100001111001000010100010",
4049 => "0010100100011010100110001",
4050 => "0010100111011010001100011",
4051 => "0101000010001101001010001",
4052 => "0101001000001100011000011",
4053 => "0011000000001100100110001",
4054 => "0100000000000100100100011",
4055 => "0011001001011000010010001",
4056 => "0011001011011000001000010",
4057 => "0001100010011110110010001",
4058 => "0001100110011110010000011",
4059 => "0110000000011000010110001",
4060 => "1000000000001000010100011",
4061 => "0000001111100100001110001",
4062 => "0011001111001100001100011",
4063 => "0000001110110000010110001",
4064 => "0100001110010000010100011",
4065 => "0010100001000111001010001",
4066 => "0011000001000011001000011",
4067 => "0101000000001000111010001",
4068 => "0101000000000100111000010",
4069 => "0100100011001000100110001",
4070 => "0101100011000100100100010",
4071 => "0100000010011000011010001",
4072 => "0111000010001100001100010",
4073 => "0100000101001100001100010",
4074 => "0000000100100010010010001",
4075 => "0000000110100010001000010",
4076 => "1000010000001010100010001",
4077 => "1000010100001010010000010",
4078 => "0001110000001010100010001",
4079 => "0001110100001010010000010",
4080 => "0011010010100100001010001",
4081 => "0011010011100100000100010",
4082 => "0000000000011000010110001",
4083 => "0010000000001000010100011",
4084 => "0111000011001100110010001",
4085 => "1000100011000110011000010",
4086 => "0111001001000110011000010",
4087 => "0000001100001100110010001",
4088 => "0001001100000100110000011",
4089 => "0001000011101010001110001",
4090 => "0001000100101010000100011",
4091 => "0010000011001100110010001",
4092 => "0010000011000110011000010",
4093 => "0011101001000110011000010",
4094 => "0110001000011000011010001",
4095 => "1001001000001100001100010",
4096 => "0110001011001100001100010",
4097 => "0000001111100000100110001",
4098 => "0100001111010000100100010",
4099 => "0011001101100100010110001",
4100 => "0011001101010010010100010",
4101 => "0000100110011110011010001",
4102 => "0011000110001010011000011",
4103 => "0101101001010010011010001",
4104 => "0111001001000110011000011",
4105 => "0001100000011110101110001",
4106 => "0100000000001010101100011",
4107 => "0111100011000111001010001",
4108 => "0111101001000110011000011",
4109 => "0011000011000111001010001",
4110 => "0011001001000110011000011",
4111 => "0100100101010100100010001",
4112 => "0111000101001010010000010",
4113 => "0100101001001010010000010",
4114 => "0010000100100000100010001",
4115 => "0010000100010000010000010",
4116 => "0110001000010000010000010",
4117 => "0011100111011000001110001",
4118 => "0011100111001100001100010",
4119 => "0010100000010010110110001",
4120 => "0100000000000110110100011",
4121 => "0101100000001100100110001",
4122 => "0110100000000100100100011",
4123 => "0011100000001100100110001",
4124 => "0100100000000100100100011",
4125 => "0100000001010100100110001",
4126 => "0100000100010100001100011",
4127 => "0000000010100100001010001",
4128 => "0000000011100100000100010",
4129 => "0101001101011100011010001",
4130 => "1000101101001110001100010",
4131 => "0101010000001110001100010",
4132 => "0000001101011100011010001",
4133 => "0000001101001110001100010",
4134 => "0011110000001110001100010",
4135 => "1010000010000111010110001",
4136 => "1010100010000011010100011",
4137 => "0000001001001010110010001",
4138 => "0000001101001010010000011",
4139 => "0110000110011000011010001",
4140 => "0110001000011000001000011",
4141 => "0000101000101000001110001",
4142 => "0000101001101000000100011",
4143 => "0010100111100110001110001",
4144 => "0010101000100110000100011",
4145 => "0000101100010010011010001",
4146 => "0000101110010010001000011",
4147 => "0011001010011100110010001",
4148 => "0011001110011100010000011",
4149 => "0010100110011101001010001",
4150 => "0010101100011100011000011",
4151 => "0101101100010010011110001",
4152 => "0111001100000110011100011",
4153 => "0000101111100100010010001",
4154 => "0000110001100100001000010",
4155 => "0101101110001100100110001",
4156 => "0101110001001100001100011",
4157 => "0000001000100100010010001",
4158 => "0000001000010010001000010",
4159 => "0100101010010010001000010",
4160 => "0001101010101000011010001",
4161 => "0110101010010100001100010",
4162 => "0001101101010100001100010",
4163 => "0000101010101000011010001",
4164 => "0000101010010100001100010",
4165 => "0101101101010100001100010",
4166 => "0000001001110000001010001",
4167 => "0000001001011000001000010",
4168 => "0000101100101000100010001",
4169 => "0000101100010100010000010",
4170 => "0101110000010100010000010",
4171 => "0101101100010010011110001",
4172 => "0111001100000110011100011",
4173 => "0010001100010010011110001",
4174 => "0011101100000110011100011",
4175 => "0110001100010000010110001",
4176 => "0110001100001000010100010",
4177 => "0010001100010000010110001",
4178 => "0100001100001000010100010",
4179 => "0110101010001000101010001",
4180 => "0110101010000100101000010",
4181 => "0000101111101000001010001",
4182 => "0101101111010100001000010",
4183 => "0100101010001100011010001",
4184 => "0100101010000110011000010",
4185 => "0000000001101010001110001",
4186 => "0011100001001110001100011",
4187 => "0011000100011010100110001",
4188 => "0011000111011010001100011",
4189 => "0011000101011000010110001",
4190 => "0101000101001000010100011",
4191 => "0101001010010100011010001",
4192 => "0101001100010100001000011",
4193 => "0011001100001010100010001",
4194 => "0011010000001010010000010",
4195 => "0110100000001100100110001",
4196 => "0111100000000100100100011",
4197 => "0001001010100100011010001",
4198 => "0100001010001100011000011",
4199 => "0101100010010010010010001",
4200 => "0101100100010010001000010",
4201 => "0000110100101010001110001",
4202 => "0100010100001110001100011",
4203 => "0000101010101100001010001",
4204 => "0000101011101100000100010",
4205 => "0000010001100100001110001",
4206 => "0000010010100100000100011",
4207 => "0110100000001100100110001",
4208 => "0111100000000100100100011",
4209 => "0010100000001100100110001",
4210 => "0011100000000100100100011",
4211 => "1001000010001101010010001",
4212 => "1010000010000101010000011",
4213 => "0000000010001101010010001",
4214 => "0001000010000101010000011",
4215 => "0101100111001100111010001",
4216 => "0111000111000110011100010",
4217 => "0101101110000110011100010",
4218 => "0000000001001000100110001",
4219 => "0001000001000100100100010",
4220 => "0110001110010010010010001",
4221 => "0110010000010010001000010",
4222 => "0000101101010010010010001",
4223 => "0000101111010010001000010",
4224 => "0011100110011110011010001",
4225 => "0011101000011110001000011",
4226 => "0100000010000111001010001",
4227 => "0100001000000110011000011",
4228 => "0011000110011000011010001",
4229 => "0110000110001100001100010",
4230 => "0011001001001100001100010",
4231 => "0001010011101000010010001",
4232 => "0001010011010100001000010",
4233 => "0110010101010100001000010",
4234 => "0111001111001100100110001",
4235 => "0111010010001100001100011",
4236 => "0001100101100100111010001",
4237 => "0001100101010010011100010",
4238 => "0110001100010010011100010",
4239 => "0111100110001001001010001",
4240 => "1000100110000100100100010",
4241 => "0111101111000100100100010",
4242 => "0010100110001001001010001",
4243 => "0010100110000100100100010",
4244 => "0011101111000100100100010",
4245 => "0101100000001100100110001",
4246 => "0110100000000100100100011",
4247 => "0011100000001100100110001",
4248 => "0100100000000100100100011",
4249 => "0101100101001100100110001",
4250 => "0110100101000100100100011",
4251 => "0100100101001100011010001",
4252 => "0110000101000110011000010",
4253 => "0010000001100000011010001",
4254 => "0110000001010000001100010",
4255 => "0010000100010000001100010",
4256 => "0100101101001100101110001",
4257 => "0101101101000100101100011",
4258 => "1000100001001100110010001",
4259 => "1010000001000110011000010",
4260 => "1000100111000110011000010",
4261 => "0000110001100100001110001",
4262 => "0000110010100100000100011",
4263 => "0011101101010100100010001",
4264 => "0011110001010100010000010",
4265 => "0011010010010100011010001",
4266 => "0011010100010100001000011",
4267 => "0100101110010010010010001",
4268 => "0100110000010010001000010",
4269 => "0000100001001100110010001",
4270 => "0000100001000110011000010",
4271 => "0010000111000110011000010",
4272 => "1001100100001010110010001",
4273 => "1001101000001010010000011",
4274 => "0000000000010000100010001",
4275 => "0010000000001000100000010",
4276 => "0001100101100110001110001",
4277 => "0001100110100110000100011",
4278 => "0000100101011000011010001",
4279 => "0000100101001100001100010",
4280 => "0011101000001100001100010",
4281 => "0001000001101010100010001",
4282 => "0100100001001110100000011",
4283 => "0010000001100000100010001",
4284 => "0010000101100000010000010",
4285 => "0011000000100100001110001",
4286 => "0011000001100100000100011",
4287 => "0010000100010100111010001",
4288 => "0010001011010100011100010",
4289 => "0111100110001000101010001",
4290 => "0111101011001000010100010",
4291 => "0001110010100100001110001",
4292 => "0100110010001100001100011",
4293 => "0100010010011000011010001",
4294 => "0110010010001000011000011",
4295 => "0001101111001100100110001",
4296 => "0011001111000110100100010",
4297 => "0111100111001100100010001",
4298 => "0111101011001100010000010",
4299 => "0001100111001100100010001",
4300 => "0001101011001100010000010",
4301 => "0010101001100100011010001",
4302 => "0111001001010010001100010",
4303 => "0010101100010010001100010",
4304 => "0000101101011000011010001",
4305 => "0000101111011000001000011",
4306 => "0111001111010100011010001",
4307 => "0111010001010100001000011",
4308 => "0000001111010100011010001",
4309 => "0000010001010100001000011",
4310 => "0111101101001100100110001",
4311 => "0111110000001100001100011",
4312 => "0001101101001100100110001",
4313 => "0001110000001100001100011",
4314 => "0100100101010000100010001",
4315 => "0100100101001000100000010",
4316 => "0000110010011000011010001",
4317 => "0000110010001100001100010",
4318 => "0011110101001100001100010",
4319 => "0110110011010100010010001",
4320 => "0110110101010100001000010",
4321 => "0000110011010100010010001",
4322 => "0000110101010100001000010",
4323 => "0011010011100100001110001",
4324 => "0011010100100100000100011",
4325 => "0100001110001000101010001",
4326 => "0100010011001000010100010",
4327 => "0000000000110000011010001",
4328 => "0000000010110000001000011",
4329 => "0000000001001100100110001",
4330 => "0000000100001100001100011",
4331 => "0010001001101000011010001",
4332 => "0111001001010100001100010",
4333 => "0010001100010100001100010",
4334 => "0000101111100110100010001",
4335 => "0000110011100110010000010",
4336 => "0111000000010100011010001",
4337 => "0111000010010100001000011",
4338 => "0000101010101010111010001",
4339 => "0100001010001110111000011",
4340 => "0101001010010000100010001",
4341 => "0101001010001000100000010",
4342 => "0011001000010100010010001",
4343 => "0101101000001010010000010",
4344 => "0101000101001000100110001",
4345 => "0101000101000100100100010",
4346 => "0011100101001100101010001",
4347 => "0100100101000100101000011",
4348 => "0111000100001000110110001",
4349 => "0111000100000100110100010",
4350 => "0011000100001000110110001",
4351 => "0100000100000100110100010",
4352 => "0100000111010010011010001",
4353 => "0101100111000110011000011",
4354 => "0001100110100000011010001",
4355 => "0001100110010000001100010",
4356 => "0101101001010000001100010",
4357 => "0010100100100000111010001",
4358 => "0110100100010000011100010",
4359 => "0010101011010000011100010",
4360 => "0000000000110000010010001",
4361 => "0000000000011000001000010",
4362 => "0110000010011000001000010",
4363 => "0100100001010010011010001",
4364 => "0110000001000110011000011",
4365 => "0010000001011100010010001",
4366 => "0101100001001110010000010",
4367 => "0101001110001110100110001",
4368 => "0101010001001110001100011",
4369 => "0100000011010000101010001",
4370 => "0100000011001000010100010",
4371 => "0110001000001000010100010",
4372 => "0011100011011000010110001",
4373 => "0101100011001000010100011",
4374 => "0100000010001000110110001",
4375 => "0101000010000100110100010",
4376 => "0101100010000111001110001",
4377 => "0110000010000011001100011",
4378 => "0011100111010010011010001",
4379 => "0101000111000110011000011",
4380 => "0010010110101000001010001",
4381 => "0010010110010100001000010",
4382 => "0000010000110000010010001",
4383 => "0000010000011000001000010",
4384 => "0110010010011000001000010",
4385 => "0011100011011000010110001",
4386 => "0101100011001000010100011",
4387 => "0000101010010000111010001",
4388 => "0000101010001000011100010",
4389 => "0010110001001000011100010",
4390 => "0101110000001100011010001",
4391 => "0101110011001100001100010",
4392 => "0011000000010101100010001",
4393 => "0011000000001010110000010",
4394 => "0101101100001010110000010",
4395 => "0011100101011100111010001",
4396 => "0111000101001110011100010",
4397 => "0011101100001110011100010",
4398 => "0011101000010100100010001",
4399 => "0011101000001010010000010",
4400 => "0110001100001010010000010",
4401 => "0100100001010010011010001",
4402 => "0110000001000110011000011",
4403 => "0000000110110000001110001",
4404 => "0110000110011000001100010",
4405 => "0011100011011000010110001",
4406 => "0101100011001000010100011",
4407 => "0000101101101100010010001",
4408 => "0000101101010110001000010",
4409 => "0110001111010110001000010",
4410 => "0100101100011000011010001",
4411 => "0100101110011000001000011",
4412 => "0000000101010010011010001",
4413 => "0000000111010010001000011",
4414 => "0000100101101110011010001",
4415 => "0000100111101110001000011",
4416 => "0000100110100110110010001",
4417 => "0000101010100110010000011",
4418 => "0100100001001101010110001",
4419 => "0100101000001100011100011",
4420 => "0001110011100100001110001",
4421 => "0100110011001100001100011",
4422 => "0100101110001100100110001",
4423 => "0101101110000100100100011",
4424 => "0100100110001000110010001",
4425 => "0101100110000100110000010",
4426 => "1000000000001100100110001",
4427 => "1001000000000100100100011",
4428 => "0001000000001100100110001",
4429 => "0010000000000100100100011",
4430 => "0110100001001001011010001",
4431 => "0111100001000100101100010",
4432 => "0110101100000100101100010",
4433 => "0000101000010000110010001",
4434 => "0000101110010000011000010",
4435 => "0111000111001110100110001",
4436 => "0111001010001110001100011",
4437 => "0001101100100100010010001",
4438 => "0001101100010010001000010",
4439 => "0110001110010010001000010",
4440 => "0110100001001001011010001",
4441 => "0111100001000100101100010",
4442 => "0110101100000100101100010",
4443 => "0011100001001001011010001",
4444 => "0011100001000100101100010",
4445 => "0100101100000100101100010",
4446 => "0010000111101000010010001",
4447 => "0111000111010100001000010",
4448 => "0010001001010100001000010",
4449 => "0100101010001100011110001",
4450 => "0110001010000110011100010",
4451 => "0011100111010100010010001",
4452 => "0011100111001010010000010",
4453 => "0000000011001000111110001",
4454 => "0000001000001000010100011",
4455 => "0111100000010000110010001",
4456 => "1001100000001000011000010",
4457 => "0111100110001000011000010",
4458 => "0000100000010000110010001",
4459 => "0000100000001000011000010",
4460 => "0010100110001000011000010",
4461 => "0111000101001101000010001",
4462 => "1000000101000101000000011",
4463 => "0010000101001101000010001",
4464 => "0011000101000101000000011",
4465 => "0111100000001101000010001",
4466 => "1000100000000101000000011",
4467 => "0001100000001101000010001",
4468 => "0010100000000101000000011",
4469 => "0000000010110000001110001",
4470 => "0000000011110000000100011",
4471 => "0011100001010100010010001",
4472 => "0011100011010100001000010",
4473 => "0000100000101110100010001",
4474 => "0000100100101110010000010",
4475 => "0000110001100110001110001",
4476 => "0000110010100110000100011",
4477 => "0011010010100100001010001",
4478 => "0011010011100100000100010",
4479 => "0000110001010010011010001",
4480 => "0000110011010010001000011",
4481 => "0111101111001100100110001",
4482 => "0111110010001100001100011",
4483 => "0001101111001100100110001",
4484 => "0001110010001100001100011",
4485 => "0010001110101000011010001",
4486 => "0010010001101000001100010",
4487 => "0000001010001100111010001",
4488 => "0000001010000110011100010",
4489 => "0001110001000110011100010",
4490 => "0011010010100100001110001",
4491 => "0011010011100100000100011",
4492 => "0010001100010010011110001",
4493 => "0011101100000110011100011",
4494 => "0011001010100100010110001",
4495 => "0110001010001100010100011",
4496 => "0000001010100100010110001",
4497 => "0011001010001100010100011",
4498 => "0001100010100100100110001",
4499 => "0100100010001100100100011",
4500 => "0010000110010100101010001",
4501 => "0010000110001010010100010",
4502 => "0100101011001010010100010",
4503 => "1010001110001000100110001",
4504 => "1010001110000100100100010",
4505 => "0000001110001000100110001",
4506 => "0001001110000100100100010",
4507 => "0101100001001001010010001",
4508 => "0110100001000100101000010",
4509 => "0101101011000100101000010",
4510 => "0011010101011000001110001",
4511 => "0110010101001100001100010",
4512 => "0101100001001001010010001",
4513 => "0110100001000100101000010",
4514 => "0101101011000100101000010",
4515 => "0000110000010100100010001",
4516 => "0000110000001010010000010",
4517 => "0011010100001010010000010",
4518 => "0101100001001001010010001",
4519 => "0110100001000100101000010",
4520 => "0101101011000100101000010",
4521 => "0000100000000111001110001",
4522 => "0001000000000011001100011",
4523 => "0101100001001001010010001",
4524 => "0110100001000100101000010",
4525 => "0101101011000100101000010",
4526 => "0000000001001100100110001",
4527 => "0001000001000100100100011",
4528 => "0001100111100110010010001",
4529 => "0001101001100110001000010",
4530 => "0011101110010010011010001",
4531 => "0011110000010010001000011",
4532 => "1000100001001110011010001",
4533 => "1000100100001110001100010",
4534 => "0010100000011100100010001",
4535 => "0010100100011100010000010",
4536 => "1000000001010000011010001",
4537 => "1000000100010000001100010",
4538 => "0000000001010000011010001",
4539 => "0000000100010000001100010",
4540 => "0011000000100100010010001",
4541 => "0111100000010010001000010",
4542 => "0011000010010010001000010",
4543 => "0000001110010010011010001",
4544 => "0000010000010010001000011",
4545 => "0001100111100100100010001",
4546 => "0100100111001100100000011",
4547 => "0001001011001100100110001",
4548 => "0010001011000100100100011",
4549 => "0101000101001100100110001",
4550 => "0110000101000100100100011",
4551 => "0101000110001001001010001",
4552 => "0101000110000100100100010",
4553 => "0110001111000100100100010",
4554 => "0101100001001001010010001",
4555 => "0110100001000100101000010",
4556 => "0101101011000100101000010",
4557 => "0100100001001001010010001",
4558 => "0100100001000100101000010",
4559 => "0101101011000100101000010",
4560 => "0010101001100100011010001",
4561 => "0111001001010010001100010",
4562 => "0010101100010010001100010",
4563 => "0011000100001100100110001",
4564 => "0100000100000100100100011",
4565 => "0101010000010000011010001",
4566 => "0101010000001000011000010",
4567 => "0000000000100100100010001",
4568 => "0000000000010010010000010",
4569 => "0100100100010010010000010",
4570 => "0011000101011100110010001",
4571 => "0110100101001110011000010",
4572 => "0011001011001110011000010",
4573 => "0010000011011110011110001",
4574 => "0100100011001010011100011",
4575 => "0111001100010100011010001",
4576 => "0111001110010100001000011",
4577 => "0000001011001000101010001",
4578 => "0000010000001000010100010",
4579 => "0000101010101100001110001",
4580 => "0000101011101100000100011",
4581 => "0100001001001100101010001",
4582 => "0101001001000100101000011",
4583 => "0110100010001100110010001",
4584 => "1000000010000110011000010",
4585 => "0110101000000110011000010",
4586 => "0101000110001001001010001",
4587 => "0101000110000100100100010",
4588 => "0110001111000100100100010",
4589 => "0011101000010101000010001",
4590 => "0110001000001010100000010",
4591 => "0011110000001010100000010",
4592 => "0100000001010000110010001",
4593 => "0100000001001000011000010",
4594 => "0110000111001000011000010",
4595 => "0011100001011000111010001",
4596 => "0110100001001100011100010",
4597 => "0011101000001100011100010",
4598 => "0001001110011000011010001",
4599 => "0001010000011000001000011",
4600 => "0101110000001100011010001",
4601 => "0101110011001100001100010",
4602 => "0011110000001100011010001",
4603 => "0011110011001100001100010",
4604 => "0110100100001000101010001",
4605 => "0110100100000100101000010",
4606 => "0000010011100110001110001",
4607 => "0000010100100110000100011",
4608 => "0110001000001100100010001",
4609 => "0110001100001100010000010",
4610 => "0100000001010001011010001",
4611 => "0100001100010000101100010",
4612 => "0110001000001100100010001",
4613 => "0110001100001100010000010",
4614 => "0011001000001100100010001",
4615 => "0011001100001100010000010",
4616 => "0111000101001100100110001",
4617 => "0111001000001100001100011",
4618 => "0000000110110000010010001",
4619 => "0000001000110000001000010",
4620 => "0111001100010100011010001",
4621 => "0111001110010100001000011",
4622 => "0000001100010100011010001",
4623 => "0000001110010100001000011",
4624 => "0010000110100110001110001",
4625 => "0010000111100110000100011",
4626 => "0000100110100110001110001",
4627 => "0000100111100110000100011",
4628 => "0010000000100000100110001",
4629 => "0010000011100000001100011",
4630 => "0000000001110000010110001",
4631 => "0100000001010000010100011",
4632 => "0001100110001100111110001",
4633 => "0001101011001100010100011",
4634 => "0100100110001100100110001",
4635 => "0101100110000100100100011",
4636 => "0000010001100100001110001",
4637 => "0000010010100100000100011",
4638 => "0011010110100100001010001",
4639 => "0011010111100100000100010",
4640 => "0001001100001100100110001",
4641 => "0001001111001100001100011",
4642 => "1001001100001100100110001",
4643 => "1001001111001100001100011",
4644 => "0000001100001100100110001",
4645 => "0000001111001100001100011",
4646 => "0101101110001000101010001",
4647 => "0101110011001000010100010",
4648 => "0100100110001101000010001",
4649 => "0100101110001100100000010",
4650 => "0011100111010100101010001",
4651 => "0011101100010100010100010",
4652 => "0000100011001100110110001",
4653 => "0001100011000100110100011",
4654 => "1001000001001100110110001",
4655 => "1001000001000110110100010",
4656 => "0010100001001100100110001",
4657 => "0011100001000100100100011",
4658 => "1001000010001100101110001",
4659 => "1001000010000110101100010",
4660 => "0000000010001100101110001",
4661 => "0001100010000110101100010",
4662 => "0100101100011110011010001",
4663 => "0100101110011110001000011",
4664 => "0001000010101000001110001",
4665 => "0001000011101000000100011",
4666 => "0101000110001000100110001",
4667 => "0101000110000100100100010",
4668 => "0010100110011000111010001",
4669 => "0010100110001100011100010",
4670 => "0101101101001100011100010",
4671 => "0100100000001100100110001",
4672 => "0101100000000100100100011",
4673 => "0011100000010010011010001",
4674 => "0101000000000110011000011",
4675 => "0101000110001100100110001",
4676 => "0110000110000100100100011",
4677 => "0010000001011001010010001",
4678 => "0010000001001100101000010",
4679 => "0101001011001100101000010",
4680 => "0011000111100100001110001",
4681 => "0011000111010010001100010",
4682 => "0000000111100100001110001",
4683 => "0100100111010010001100010",
4684 => "0001110100100100001110001",
4685 => "0100110100001100001100011",
4686 => "0100100110001100100110001",
4687 => "0101100110000100100100011",
4688 => "0011000010011000111110001",
4689 => "0101000010001000111100011",
4690 => "0001000011100100001110001",
4691 => "0001000100100100000100011",
4692 => "1001100100001001001010001",
4693 => "1010100100000100100100010",
4694 => "1001101101000100100100010",
4695 => "0000000001100110001110001",
4696 => "0000000010100110000100011",
4697 => "0010100000011110010010001",
4698 => "0010100010011110001000010",
4699 => "0010100010011100010110001",
4700 => "0110000010001110010100010",
4701 => "0000100010101100111010001",
4702 => "0000100010010110111000010",
4703 => "0100001111001100100110001",
4704 => "0101001111000100100100011",
4705 => "0011010001100100001110001",
4706 => "0011010010100100000100011",
4707 => "0100100110000111001010001",
4708 => "0100101100000110011000011",
4709 => "0001000000101000001110001",
4710 => "0001000001101000000100011",
4711 => "0010100100001010110010001",
4712 => "0010101000001010010000011",
4713 => "0100000110011000010110001",
4714 => "0110000110001000010100011",
4715 => "0100101100001100110010001",
4716 => "0100101100000110011000010",
4717 => "0110010010000110011000010",
4718 => "0111001110010000101010001",
4719 => "1001001110001000010100010",
4720 => "0111010011001000010100010",
4721 => "0001001110010000101010001",
4722 => "0001001110001000010100010",
4723 => "0011010011001000010100010",
4724 => "0101010010011000011010001",
4725 => "1000010010001100001100010",
4726 => "0101010101001100001100010",
4727 => "0000100011001100100110001",
4728 => "0000100110001100001100011",
4729 => "0101100011000111010010001",
4730 => "0110000011000011010000011",
4731 => "0010000110011100011010001",
4732 => "0010000110001110001100010",
4733 => "0101101001001110001100010",
4734 => "0011000101011000110110001",
4735 => "0101000101001000110100011",
4736 => "0010100100001000111110001",
4737 => "0010101001001000010100011",
4738 => "0100110000011110010010001",
4739 => "0111010000001010010000011",
4740 => "0011101000001100111010001",
4741 => "0011101000000110011100010",
4742 => "0101001111000110011100010",
4743 => "0011100110010100011010001",
4744 => "0011101000010100001000011",
4745 => "0001000101100100001110001",
4746 => "0001000110100100000100011",
4747 => "0010100001011110100010001",
4748 => "0010100101011110010000010",
4749 => "0011100001010001001010001",
4750 => "0011101010010000100100010",
4751 => "0000001010110000001110001",
4752 => "0000001011110000000100011",
4753 => "0000000010001100110110001",
4754 => "0001000010000100110100011",
4755 => "1000000000010000101010001",
4756 => "1010000000001000010100010",
4757 => "1000000101001000010100010",
4758 => "0010100001010100100110001",
4759 => "0010100100010100001100011",
4760 => "0010100110100100001110001",
4761 => "0010100111100100000100011",
4762 => "0000000001110000001110001",
4763 => "0000000010110000000100011",
4764 => "0101100100001100101110001",
4765 => "0110100100000100101100011",
4766 => "0000000000010000101010001",
4767 => "0000000000001000010100010",
4768 => "0010000101001000010100010",
4769 => "0010010000100100001110001",
4770 => "0010010001100100000100011",
4771 => "0001010000100100001110001",
4772 => "0001010001100100000100011",
4773 => "0001100000100100101010001",
4774 => "0110000000010010010100010",
4775 => "0001100101010010010100010",
4776 => "0001000011101001010110001",
4777 => "0110000011010101010100010",
4778 => "0011000111011100001110001",
4779 => "0011000111001110001100010",
4780 => "0000001001011000011010001",
4781 => "0000001001001100001100010",
4782 => "0011001100001100001100010",
4783 => "0001101110101010010010001",
4784 => "0101001110001110010000011",
4785 => "0000001110101010010010001",
4786 => "0011101110001110010000011",
4787 => "0010110101100100001110001",
4788 => "0101110101001100001100011",
4789 => "0000110101100100001110001",
4790 => "0011110101001100001100011",
4791 => "1001100100001001001010001",
4792 => "1010100100000100100100010",
4793 => "1001101101000100100100010",
4794 => "0001100111100100001110001",
4795 => "0001101000100100000100011",
4796 => "1001100100001001001010001",
4797 => "1010100100000100100100010",
4798 => "1001101101000100100100010",
4799 => "0011101111010100011010001",
4800 => "0011110001010100001000011",
4801 => "0100101101010110100110001",
4802 => "0100110000010110001100011",
4803 => "0000000110001000101010001",
4804 => "0000001011001000010100010",
4805 => "0111110000010010011010001",
4806 => "0111110010010010001000011",
4807 => "0000100101001001001010001",
4808 => "0000100101000100100100010",
4809 => "0001101110000100100100010",
4810 => "0100101000010000101010001",
4811 => "0110101000001000010100010",
4812 => "0100101101001000010100010",
4813 => "0011101000010000101010001",
4814 => "0011101000001000010100010",
4815 => "0101101101001000010100010",
4816 => "0100101000011000010110001",
4817 => "0110101000001000010100011",
4818 => "0011101000010010011110001",
4819 => "0101001000000110011100011",
4820 => "0100101000011000010110001",
4821 => "0110101000001000010100011",
4822 => "0011100110010010011110001",
4823 => "0101000110000110011100011",
4824 => "0100101000011000010110001",
4825 => "0110101000001000010100011",
4826 => "0101000101001001001010001",
4827 => "0101001011001000011000011",
4828 => "0010100101011100110010001",
4829 => "0010101011011100011000010",
4830 => "0000000001010110010010001",
4831 => "0000000011010110001000010",
4832 => "0100101010001100101010001",
4833 => "0101101010000100101000011",
4834 => "0001010001010110011010001",
4835 => "0001010011010110001000011",
4836 => "0111110000010010011010001",
4837 => "0111110010010010001000011",
4838 => "0000101010100100001010001",
4839 => "0000101011100100000100010",
4840 => "0011000100011000110110001",
4841 => "0101000100001000110100011",
4842 => "0000010010100100001110001",
4843 => "0000010011100100000100011",
4844 => "0011010010100100001110001",
4845 => "0011010011100100000100011",
4846 => "0000010000010010011010001",
4847 => "0000010010010010001000011",
4848 => "0110101111010010011010001",
4849 => "0110110001010010001000011",
4850 => "0001001111010010011010001",
4851 => "0001010001010010001000011",
4852 => "0110100001001101000010001",
4853 => "0110100001000111000000010",
4854 => "0010100001001101000010001",
4855 => "0100000001000111000000010",
4856 => "0101100101001100101010001",
4857 => "0110100101000100101000011",
4858 => "0011100101001100101010001",
4859 => "0100100101000100101000011",
4860 => "0101000000001101100010001",
4861 => "0110000000000101100000011",
4862 => "0001100100001001010010001",
4863 => "0001100100000100101000010",
4864 => "0010101110000100101000010",
4865 => "0111000000001100100110001",
4866 => "1000000000000100100100011",
4867 => "0010000000001100100110001",
4868 => "0011000000000100100100011",
4869 => "0010000101100100010110001",
4870 => "0101000101001100010100011",
4871 => "0010100110001100100110001",
4872 => "0011100110000100100100011",
4873 => "0011100010011110100010001",
4874 => "0110000010001010100000011",
4875 => "0001000010011110100010001",
4876 => "0011100010001010100000011",
4877 => "0101000000001000100110001",
4878 => "0101000000000100100100010",
4879 => "0001100100001100110010001",
4880 => "0001100100000110011000010",
4881 => "0011001010000110011000010",
4882 => "1000000000010001001010001",
4883 => "1000000000001001001000010",
4884 => "0000000000010001001010001",
4885 => "0010000000001001001000010",
4886 => "0000000111110000011010001",
4887 => "0000001001110000001000011",
4888 => "0010000111011100001110001",
4889 => "0101100111001110001100010",
4890 => "0101001000010000111110001",
4891 => "0101001000001000111100010",
4892 => "0011100000010100111010001",
4893 => "0110000000001010111000010",
4894 => "0110101010010000101010001",
4895 => "1000101010001000010100010",
4896 => "0110101111001000010100010",
4897 => "0001100000001000100110001",
4898 => "0010100000000100100100010",
4899 => "1000000001001100100010001",
4900 => "1000000001000110100000010",
4901 => "0001000001001100100010001",
4902 => "0010100001000110100000010",
4903 => "0001100110100100110010001",
4904 => "0001101010100100010000011",
4905 => "0010001100100000010010001",
4906 => "0010001110100000001000010",
4907 => "0010001001100000111110001",
4908 => "0010001110100000010100011",
4909 => "0001101010010000101010001",
4910 => "0001101010001000010100010",
4911 => "0011101111001000010100010",
4912 => "0100010010100000011010001",
4913 => "1000010010010000001100010",
4914 => "0100010101010000001100010",
4915 => "0001010000011000010110001",
4916 => "0011010000001000010100011",
4917 => "0111001110010010010010001",
4918 => "0111010000010010001000010",
4919 => "0011101110010010011010001",
4920 => "0011110000010010001000011",
4921 => "0010001010100000110010001",
4922 => "0010001110100000010000011",
4923 => "0000001101100110011010001",
4924 => "0000001111100110001000011",
4925 => "0101001101010010011010001",
4926 => "0101001111010010001000011",
4927 => "0010100000000111011110001",
4928 => "0011000000000011011100011",
4929 => "0000001000110000011010001",
4930 => "0000001010110000001000011",
4931 => "0000000101001010110010001",
4932 => "0000001001001010010000011",
4933 => "0001100000100111001010001",
4934 => "0001101001100110100100010",
4935 => "0100101011001100110010001",
4936 => "0100101011000110011000010",
4937 => "0110010001000110011000010",
4938 => "0000000101110000100010001",
4939 => "0110000101011000010000010",
4940 => "0000001001011000010000010",
4941 => "0011010010010010010010001",
4942 => "0011010100010010001000010",
4943 => "0100001000010100011010001",
4944 => "0100001010010100001000011",
4945 => "0001000111101000001110001",
4946 => "0001001000101000000100011",
4947 => "0110000000001111010010001",
4948 => "0110001010001110101000010",
4949 => "0010100000001111010010001",
4950 => "0010101010001110101000010",
4951 => "0111000010000101001010001",
4952 => "0111001011000100100100010",
4953 => "0010101000010100110010001",
4954 => "0101001000001010110000010",
4955 => "0011001001011000100010001",
4956 => "0110001001001100010000010",
4957 => "0011001101001100010000010",
4958 => "0011100111000110111010001",
4959 => "0011101110000110011100010",
4960 => "0101100010011001000010001",
4961 => "1000100010001100100000010",
4962 => "0101101010001100100000010",
4963 => "0011100000001100100110001",
4964 => "0100100000000100100100011",
4965 => "0110101110010010010010001",
4966 => "0110110000010010001000010",
4967 => "0000001100101100010010001",
4968 => "0000001100010110001000010",
4969 => "0101101110010110001000010",
4970 => "0000101100101100011010001",
4971 => "0110001100010110001100010",
4972 => "0000101111010110001100010",
4973 => "0011000110010010011010001",
4974 => "0100100110000110011000011",
4975 => "0101000000001000100110001",
4976 => "0101000000000100100100010",
4977 => "0001101000100100011110001",
4978 => "0100101000001100011100011",
4979 => "0000000110110000011010001",
4980 => "0000001000110000001000011",
4981 => "0000001011110000101010001",
4982 => "0100001011010000101000011",
4983 => "0001100011100101010110001",
4984 => "0100100011001101010100011",
4985 => "0011101100001000101010001",
4986 => "0100101100000100101000010",
4987 => "0101010000010100100010001",
4988 => "0111110000001010010000010",
4989 => "0101010100001010010000010",
4990 => "0100000110001100100110001",
4991 => "0101000110000100100100011",
4992 => "0110001010001100110010001",
4993 => "0111101010000110011000010",
4994 => "0110010000000110011000010",
4995 => "0011001010001100110010001",
4996 => "0011001010000110011000010",
4997 => "0100110000000110011000010",
4998 => "1000001100001100110010001",
4999 => "1001101100000110011000010",
5000 => "1000010010000110011000010",
5001 => "0001001100001100110010001",
5002 => "0001001100000110011000010",
5003 => "0010110010000110011000010",
5004 => "0101001111001100100110001",
5005 => "0110001111000100100100011",
5006 => "0100001111001100100110001",
5007 => "0101001111000100100100011",
5008 => "0111010100010100010010001",
5009 => "0111010100001010010000010",
5010 => "0000010100010100010010001",
5011 => "0010110100001010010000010",
5012 => "0101110001010010011010001",
5013 => "0101110011010010001000011",
5014 => "0001100010011100010010001",
5015 => "0001100100011100001000010",
5016 => "0101000001010100010010001",
5017 => "0101000011010100001000010",
5018 => "0000001111010100010010001",
5019 => "0010101111001010010000010",
5020 => "1001100010000111001110001",
5021 => "1010000010000011001100011",
5022 => "0010001100010010100010001",
5023 => "0011101100000110100000011",
5024 => "0010000111001010110010001",
5025 => "0010001011001010010000011",
5026 => "0000000001110000001110001",
5027 => "0100000001010000001100011",
5028 => "0011001000011000010010001",
5029 => "0011001010011000001000010",
5030 => "1001100011001000101010001",
5031 => "1001100011000100101000010",
5032 => "0000000110010010011010001",
5033 => "0001100110000110011000011",
5034 => "1001000000001101011010001",
5035 => "1010000000000101011000011",
5036 => "0000000000001101011010001",
5037 => "0001000000000101011000011",
5038 => "0010101111100110001110001",
5039 => "0010110000100110000100011",
5040 => "0101000111001000111110001",
5041 => "0101001100001000010100011",
5042 => "0100100110001100100110001",
5043 => "0101100110000100100100011",
5044 => "0000010101100100001110001",
5045 => "0000010110100100000100011",
5046 => "0011100011010100111110001",
5047 => "0011101000010100010100011",
5048 => "0000100111100100001110001",
5049 => "0000101000100100000100011",
5050 => "0100000010010010011010001",
5051 => "0101100010000110011000011",
5052 => "0000001010110000111010001",
5053 => "0000010001110000011100010",
5054 => "0110101001010000101010001",
5055 => "1000101001001000010100010",
5056 => "0110101110001000010100010",
5057 => "0101000101001000100110001",
5058 => "0110000101000100100100010",
5059 => "0110101001010000101010001",
5060 => "1000101001001000010100010",
5061 => "0110101110001000010100010",
5062 => "0011101011010100101010001",
5063 => "0011101011001010010100010",
5064 => "0110010000001010010100010",
5065 => "0010001101100100010010001",
5066 => "0110101101010010001000010",
5067 => "0010001111010010001000010",
5068 => "0000000000100110001010001",
5069 => "0000000001100110000100010",
5070 => "0000010010110000011010001",
5071 => "0100010010010000011000011",
5072 => "0011000100010001000010001",
5073 => "0011001100010000100000010",
5074 => "0011101000010100010010001",
5075 => "0011101010010100001000010",
5076 => "0000000011001100100110001",
5077 => "0000000110001100001100011",
5078 => "0110101111001110100110001",
5079 => "0110110010001110001100011",
5080 => "0001110010011000011010001",
5081 => "0001110010001100001100010",
5082 => "0100110101001100001100010",
5083 => "0110001110001100100110001",
5084 => "0110010001001100001100011",
5085 => "0001001111011110100010001",
5086 => "0001010011011110010000010",
5087 => "0100100110001101000010001",
5088 => "0100101110001100100000010",
5089 => "0011000110001110110010001",
5090 => "0011001010001110010000011",
5091 => "0111000110001100100110001",
5092 => "0111001001001100001100011",
5093 => "0010101110001100100110001",
5094 => "0010110001001100001100011",
5095 => "0101001000001100100110001",
5096 => "0110001000000100100100011",
5097 => "0011000110001001001010001",
5098 => "0011000110000100100100010",
5099 => "0100001111000100100100010",
5100 => "0111001001001100110010001",
5101 => "1000101001000110011000010",
5102 => "0111001111000110011000010",
5103 => "0010001001001100110010001",
5104 => "0010001001000110011000010",
5105 => "0011101111000110011000010",
5106 => "0111001111010010011010001",
5107 => "0111010001010010001000011",
5108 => "0000010100100100010010001",
5109 => "0000010100010010001000010",
5110 => "0100110110010010001000010",
5111 => "0110110010010010011010001",
5112 => "0110110100010010001000011",
5113 => "0001010010010010011010001",
5114 => "0001010100010010001000011",
5115 => "0011010000100100001110001",
5116 => "0011010001100100000100011",
5117 => "0000010000100100001110001",
5118 => "0000010001100100000100011",
5119 => "1001100010001001011010001",
5120 => "1010100010000100101100010",
5121 => "1001101101000100101100010",
5122 => "0000100010001001011010001",
5123 => "0000100010000100101100010",
5124 => "0001101101000100101100010",
5125 => "0111100000000101100010001",
5126 => "0111100000000011100000010",
5127 => "0001110100100000010010001",
5128 => "0101110100010000010000010",
5129 => "0101100110001001001010001",
5130 => "0110100110000100100100010",
5131 => "0101101111000100100100010",
5132 => "0011101001010100111010001",
5133 => "0011101001001010011100010",
5134 => "0110010000001010011100010",
5135 => "0111000110001100100110001",
5136 => "0111001001001100001100011",
5137 => "0001100110001110100110001",
5138 => "0001101001001110001100011",
5139 => "1010000100001001010010001",
5140 => "1011000100000100101000010",
5141 => "1010001110000100101000010",
5142 => "0011100110001100100110001",
5143 => "0011101001001100001100011",
5144 => "0011100000010100111010001",
5145 => "0110000000001010011100010",
5146 => "0011100111001010011100010",
5147 => "0001000001100100011010001",
5148 => "0101100001010010011000010",
5149 => "0111100000000101100010001",
5150 => "0111100000000011100000010",
5151 => "0011100000000101100010001",
5152 => "0100000000000011100000010",
5153 => "0110101100001100011110001",
5154 => "0110101100000110011100010",
5155 => "0010101100001100011110001",
5156 => "0100001100000110011100010",
5157 => "0001100101100101001110001",
5158 => "0100100101001101001100011",
5159 => "0010100110010010011010001",
5160 => "0100000110000110011000011",
5161 => "0100100101010010011010001",
5162 => "0110000101000110011000011",
5163 => "0001110000010100100010001",
5164 => "0001110000001010010000010",
5165 => "0100010100001010010000010",
5166 => "1001101000001010111110001",
5167 => "1001101101001010010100011",
5168 => "0000001000001010111110001",
5169 => "0000001101001010010100011",
5170 => "1010000100001001010010001",
5171 => "1011000100000100101000010",
5172 => "1010001110000100101000010",
5173 => "0000000100001001010010001",
5174 => "0000000100000100101000010",
5175 => "0001001110000100101000010",
5176 => "0011100111010100010010001",
5177 => "0011100111001010010000010",
5178 => "0010010011011100010010001",
5179 => "0101110011001110010000010",
5180 => "0101001011011000001110001",
5181 => "0101001011001100001100010",
5182 => "0000000001110000001110001",
5183 => "0000000010110000000100011",
5184 => "0011100010011101010010001",
5185 => "0111000010001110101000010",
5186 => "0011101100001110101000010",
5187 => "0000001101001100100110001",
5188 => "0001001101000100100100011",
5189 => "0110100000001001001110001",
5190 => "0110100000000101001100010",
5191 => "0000101011011100001110001",
5192 => "0100001011001110001100010",
5193 => "0011100001100001010010001",
5194 => "0111100001010000101000010",
5195 => "0011101011010000101000010",
5196 => "0000001010101010100110001",
5197 => "0011101010001110100100011",
5198 => "0011010011011110010110001",
5199 => "0101110011001010010100011",
5200 => "0100001010001100011010001",
5201 => "0101101010000110011000010",
5202 => "0011100001100001010010001",
5203 => "0111100001010000101000010",
5204 => "0011101011010000101000010",
5205 => "0000100001100001010010001",
5206 => "0000100001010000101000010",
5207 => "0100101011010000101000010",
5208 => "1000000100000110110010001",
5209 => "1000001010000110011000010",
5210 => "0010100100000110110010001",
5211 => "0010101010000110011000010",
5212 => "0011100110010100100010001",
5213 => "0110000110001010010000010",
5214 => "0011101010001010010000010",
5215 => "0010001001001100011010001",
5216 => "0010001100001100001100010",
5217 => "0011000101011000010010001",
5218 => "0011000111011000001000010",
5219 => "0100100010001010111110001",
5220 => "0100100111001010010100011",
5221 => "0111100000010010011010001",
5222 => "0111100010010010001000011",
5223 => "0011000000010110101010001",
5224 => "0011000101010110010100010",
5225 => "0110000111001000110010001",
5226 => "0110001101001000011000010",
5227 => "0011100010010010010010001",
5228 => "0011100100010010001000010",
5229 => "0011000000011010011010001",
5230 => "0011000010011010001000011",
5231 => "0101000110001001001010001",
5232 => "0101000110000100100100010",
5233 => "0110001111000100100100010",
5234 => "0101001000001100100110001",
5235 => "0110001000000100100100011",
5236 => "0001110010010100011010001",
5237 => "0001110100010100001000011",
5238 => "0010001110101000001110001",
5239 => "0010001111101000000100011",
5240 => "0001001111010010011010001",
5241 => "0001010001010010001000011",
5242 => "0110100000001001001110001",
5243 => "0110100000000101001100010",
5244 => "0011100000001001001110001",
5245 => "0100100000000101001100010",
5246 => "0000100100101100001010001",
5247 => "0000100101101100000100010",
5248 => "0000000000010010011010001",
5249 => "0000000010010010001000011",
5250 => "0000000000110001001010001",
5251 => "0000001001110000100100010",
5252 => "0001100010100000100010001",
5253 => "0001100110100000010000010",
5254 => "0001100110100100011010001",
5255 => "0001101000100100001000011",
5256 => "0001100001001100101010001",
5257 => "0010100001000100101000011",
5258 => "0110100000010010011010001",
5259 => "1000000000000110011000011",
5260 => "0001000000010010011010001",
5261 => "0010100000000110011000011",
5262 => "0101000010001000111110001",
5263 => "0101000111001000010100011",
5264 => "0011000000001110101010001",
5265 => "0011000101001110010100010",
5266 => "0001000010101000010010001",
5267 => "0110000010010100001000010",
5268 => "0001000100010100001000010",
5269 => "0001001011100110001110001",
5270 => "0001001100100110000100011",
5271 => "0101001000001100100110001",
5272 => "0110001000000100100100011",
5273 => "0100001000001100100110001",
5274 => "0101001000000100100100011",
5275 => "0110101000001000100110001",
5276 => "0110101000000100100100010",
5277 => "0001101011010010100110001",
5278 => "0011001011000110100100011",
5279 => "0001101001100100010110001",
5280 => "0100101001001100010100011",
5281 => "0001000100000101010010001",
5282 => "0001001110000100101000010",
5283 => "0111010001010000011010001",
5284 => "0111010100010000001100010",
5285 => "0001110101100100001010001",
5286 => "0001110110100100000100010",
5287 => "0010100100011110011010001",
5288 => "0101000100001010011000011",
5289 => "0001001111011000011010001",
5290 => "0001010001011000001000011",
5291 => "1000101000001100100110001",
5292 => "1000101011001100001100011",
5293 => "0001001100101000010010001",
5294 => "0001001100010100001000010",
5295 => "0110001110010100001000010",
5296 => "0000010001110000011010001",
5297 => "0000010011110000001000011",
5298 => "0011110000010010010010001",
5299 => "0011110010010010001000010",
5300 => "0111100001001001011010001",
5301 => "1000100001000100101100010",
5302 => "0111101100000100101100010",
5303 => "0010100001001001011010001",
5304 => "0010100001000100101100010",
5305 => "0011101100000100101100010",
5306 => "0101101101010000100110001",
5307 => "0101110000010000001100011",
5308 => "0011000001001100100110001",
5309 => "0100000001000100100100011",
5310 => "0101100100000111001010001",
5311 => "0101101010000110011000011",
5312 => "0010101000011000011010001",
5313 => "0010101000001100001100010",
5314 => "0101101011001100001100010",
5315 => "0111100111001010100010001",
5316 => "0111101011001010010000010",
5317 => "0010000111001010100010001",
5318 => "0010001011001010010000010",
5319 => "0110000110001100110010001",
5320 => "0111100110000110011000010",
5321 => "0110001100000110011000010",
5322 => "0011000110001100110010001",
5323 => "0011000110000110011000010",
5324 => "0100101100000110011000010",
5325 => "0010101001011100100010001",
5326 => "0110001001001110010000010",
5327 => "0010101101001110010000010",
5328 => "0100100001000110111010001",
5329 => "0100101000000110011100010",
5330 => "0110000110001100110010001",
5331 => "0110001010001100010000011",
5332 => "0010000101001001001010001",
5333 => "0010000101000100100100010",
5334 => "0011001110000100100100010",
5335 => "0010000110100001001010001",
5336 => "0010001100100000011000011",
5337 => "0010100100001111010010001",
5338 => "0010101110001110101000010",
5339 => "0111001000010000110010001",
5340 => "0111001110010000011000010",
5341 => "0100101010001100111010001",
5342 => "0100101010000110011100010",
5343 => "0110010001000110011100010",
5344 => "0100100101010010011010001",
5345 => "0110000101000110011000011",
5346 => "0100100100000111001010001",
5347 => "0101000100000011001000011",
5348 => "0000100100101100111010001",
5349 => "0110000100010110011100010",
5350 => "0000101011010110011100010",
5351 => "0001000111100100001010001",
5352 => "0001001000100100000100010",
5353 => "0110000110001100110010001",
5354 => "0110001010001100010000011",
5355 => "0011000101010010011110001",
5356 => "0100100101000110011100011",
5357 => "0110000111001000110010001",
5358 => "0110001101001000011000010",
5359 => "0100000111001000110010001",
5360 => "0100001101001000011000010",
5361 => "0011100010010101011010001",
5362 => "0011101101010100101100010",
5363 => "0000000001000111010010001",
5364 => "0000100001000011010000011",
5365 => "0010001101100100010010001",
5366 => "0110101101010010001000010",
5367 => "0010001111010010001000010",
5368 => "0001001101100100010010001",
5369 => "0001001101010010001000010",
5370 => "0101101111010010001000010",
5371 => "0111101111010010011010001",
5372 => "0111110001010010001000011",
5373 => "0000001111010010011010001",
5374 => "0000010001010010001000011",
5375 => "0011000000100101100010001",
5376 => "0111100000010010110000010",
5377 => "0011001100010010110000010",
5378 => "0011000110001100110010001",
5379 => "0011001010001100010000011",
5380 => "0100000111010100010010001",
5381 => "0100001001010100001000010",
5382 => "0000101001100100011010001",
5383 => "0000101001010010001100010",
5384 => "0101001100010010001100010",
5385 => "0011000110100100001110001",
5386 => "0011000111100100000100011",
5387 => "0011100111010010100010001",
5388 => "0101000111000110100000011",
5389 => "0101001100001100110010001",
5390 => "0110001100000100110000011",
5391 => "0001101110100100001110001",
5392 => "0001101111100100000100011",
5393 => "0111110001010010011110001",
5394 => "1001010001000110011100011",
5395 => "0000101100010100011010001",
5396 => "0000101110010100001000011",
5397 => "0111110001010010011110001",
5398 => "1001010001000110011100011",
5399 => "0101000011000111001110001",
5400 => "0101100011000011001100011",
5401 => "0111110001010010011110001",
5402 => "1001010001000110011100011",
5403 => "0011000001010110100110001",
5404 => "0011000100010110001100011",
5405 => "0111110001010010011110001",
5406 => "1001010001000110011100011",
5407 => "0011000101010110011010001",
5408 => "0011001000010110001100010",
5409 => "1000000111010000010110001",
5410 => "1000000111001000010100010",
5411 => "0001000100101001001110001",
5412 => "0110000100010101001100010",
5413 => "0001000001101010011010001",
5414 => "0100100001001110011000011",
5415 => "0011000101011000111010001",
5416 => "0011000101001100011100010",
5417 => "0110001100001100011100010",
5418 => "0100100000001100100110001",
5419 => "0101100000000100100100011",
5420 => "0001001011010000010110001",
5421 => "0011001011001000010100010",
5422 => "1000000111010000010110001",
5423 => "1000000111001000010100010",
5424 => "0000000111010000010110001",
5425 => "0010000111001000010100010",
5426 => "0111110001010010011110001",
5427 => "1001010001000110011100011",
5428 => "0100000110010000101010001",
5429 => "0100000110001000010100010",
5430 => "0110001011001000010100010",
5431 => "0111101111010010100110001",
5432 => "1001001111000110100100011",
5433 => "0000001111010010100110001",
5434 => "0001101111000110100100011",
5435 => "0110001010010010011110001",
5436 => "0111101010000110011100011",
5437 => "0001101010010010011110001",
5438 => "0011001010000110011100011",
5439 => "0110101111010100100010001",
5440 => "1001001111001010010000010",
5441 => "0110110011001010010000010",
5442 => "0000000001001100110010001",
5443 => "0000000001000110011000010",
5444 => "0001100111000110011000010",
5445 => "0101000000001100110010001",
5446 => "0110100000000110011000010",
5447 => "0101000110000110011000010",
5448 => "0011100000010100110010001",
5449 => "0011100000001010011000010",
5450 => "0110000110001010011000010",
5451 => "0010000001100000100010001",
5452 => "0010000001010000100000010",
5453 => "0000010101100110001110001",
5454 => "0000010110100110000100011",
5455 => "0011001001100100010010001",
5456 => "0111101001010010001000010",
5457 => "0011001011010010001000010",
5458 => "0001100100010010011010001",
5459 => "0001100110010010001000011",
5460 => "0100100001001100111110001",
5461 => "0100100110001100010100011",
5462 => "0010101001001100011010001",
5463 => "0100001001000110011000010",
5464 => "0010100001011100100110001",
5465 => "0010100100011100001100011",
5466 => "0001100000010001010010001",
5467 => "0001100000001000101000010",
5468 => "0011101010001000101000010",
5469 => "0010100000001110100110001",
5470 => "0010100011001110001100011",
5471 => "0011000110011000010110001",
5472 => "0101000110001000010100011",
5473 => "0000000001010000111010001",
5474 => "0010000001001000111000010",
5475 => "0001001100101100010010001",
5476 => "0001001110101100001000010",
5477 => "0100010001001100011010001",
5478 => "0100010100001100001100010",
5479 => "1001000001001100011110001",
5480 => "1001000001000110011100010",
5481 => "0000000000001100011010001",
5482 => "0001100000000110011000010",
5483 => "0010000110100011001010001",
5484 => "0010001100100010011000011",
5485 => "0011000000011000011010001",
5486 => "0011000000001100001100010",
5487 => "0110000011001100001100010",
5488 => "0010000111100100010010001",
5489 => "0110100111010010001000010",
5490 => "0010001001010010001000010",
5491 => "0010001100010100011010001",
5492 => "0010001110010100001000011",
5493 => "0011101001010100110010001",
5494 => "0110001001001010011000010",
5495 => "0011101111001010011000010",
5496 => "0000000001110000001110001",
5497 => "0100000001010000001100011",
5498 => "0110101011001100011010001",
5499 => "0110101011000110011000010",
5500 => "0010101011001100011010001",
5501 => "0100001011000110011000010",
5502 => "0001101010100110001110001",
5503 => "0001101011100110000100011",
5504 => "0000000010001100100110001",
5505 => "0000000101001100001100011",
5506 => "0111010000010100011010001",
5507 => "0111010010010100001000011",
5508 => "0000010000010100011010001",
5509 => "0000010010010100001000011",
5510 => "0111001101010010011010001",
5511 => "0111001111010010001000011",
5512 => "0000010000100100001110001",
5513 => "0000010001100100000100011",
5514 => "0011010000100100001110001",
5515 => "0011010001100100000100011",
5516 => "0000010010010010011010001",
5517 => "0000010100010010001000011",
5518 => "0111001101010010011010001",
5519 => "0111001111010010001000011",
5520 => "0011000010001100100110001",
5521 => "0100000010000100100100011",
5522 => "0111101000001000110010001",
5523 => "0111101000000100110000010",
5524 => "0100001101010000100010001",
5525 => "0100010001010000010000010",
5526 => "0010010100100100001110001",
5527 => "0101010100001100001100011",
5528 => "0010101000001000110010001",
5529 => "0011101000000100110000010",
5530 => "0011100111011000001110001",
5531 => "0011100111001100001100010",
5532 => "0101000110001000100110001",
5533 => "0110000110000100100100010",
5534 => "0010110100100100001110001",
5535 => "0101110100001100001100011",
5536 => "0000110100100100001110001",
5537 => "0011110100001100001100011",
5538 => "1001000001001101010010001",
5539 => "1010100001000110101000010",
5540 => "1001001011000110101000010",
5541 => "0000000001001101010010001",
5542 => "0000000001000110101000010",
5543 => "0001101011000110101000010",
5544 => "0110100011001001001010001",
5545 => "0111100011000100100100010",
5546 => "0110101100000100100100010",
5547 => "0000000010001100110010001",
5548 => "0000000110001100010000011",
5549 => "0110001001011000011010001",
5550 => "1001001001001100001100010",
5551 => "0110001100001100001100010",
5552 => "0011100011001001001010001",
5553 => "0011100011000100100100010",
5554 => "0100101100000100100100010",
5555 => "0111000000001100100110001",
5556 => "1000000000000100100100011",
5557 => "0000001001011000011010001",
5558 => "0000001001001100001100010",
5559 => "0011001100001100001100010",
5560 => "0111000100010001010010001",
5561 => "1001000100001000101000010",
5562 => "0111001110001000101000010",
5563 => "0001000100010001010010001",
5564 => "0001000100001000101000010",
5565 => "0011001110001000101000010",
5566 => "0111001101010010011010001",
5567 => "0111001111010010001000011",
5568 => "0000101101010010011010001",
5569 => "0000101111010010001000011",
5570 => "0001101111100100001110001",
5571 => "0100101111001100001100011",
5572 => "0010101101010010011010001",
5573 => "0010101111010010001000011",
5574 => "0010100000100100001110001",
5575 => "0010100001100100000100011",
5576 => "0100000010001100011110001",
5577 => "0101100010000110011100010",
5578 => "0100100001010010011010001",
5579 => "0110000001000110011000011",
5580 => "0011000001010010011010001",
5581 => "0100100001000110011000011",
5582 => "0010100110011100011010001",
5583 => "0110000110001110001100010",
5584 => "0010101001001110001100010",
5585 => "0100000010001100110110001",
5586 => "0101000010000100110100011",
5587 => "0011001011011000011010001",
5588 => "0110001011001100001100010",
5589 => "0011001110001100001100010",
5590 => "0001100001100100111110001",
5591 => "0100100001001100111100011",
5592 => "0110100000001100011110001",
5593 => "0110100000000110011100010",
5594 => "0001100011100000011010001",
5595 => "0001100110100000001100010",
5596 => "0110000001000110110010001",
5597 => "0110000111000110011000010",
5598 => "0011100111001100100110001",
5599 => "0100100111000100100100011",
5600 => "0110100000001001100010001",
5601 => "0110100000000101100000010",
5602 => "0011100000001001100010001",
5603 => "0100100000000101100000010",
5604 => "0101101001001010110010001",
5605 => "0101101101001010010000011",
5606 => "0011101111010010011010001",
5607 => "0011110001010010001000011",
5608 => "0010100111100100011010001",
5609 => "0010101001100100001000011",
5610 => "0100001001001010110010001",
5611 => "0100001101001010010000011",
5612 => "0010010001100010011010001",
5613 => "0010010011100010001000011",
5614 => "0000000011100100111010001",
5615 => "0000000011010010011100010",
5616 => "0100101010010010011100010",
5617 => "0000000001110000001010001",
5618 => "0000000010110000000100010",
5619 => "0000001111100100001110001",
5620 => "0000010000100100000100011",
5621 => "0100100000001100100110001",
5622 => "0101100000000100100100011",
5623 => "0001100011011100110010001",
5624 => "0001101001011100011000010",
5625 => "0110000001000110110010001",
5626 => "0110000111000110011000010",
5627 => "0100000000001100100110001",
5628 => "0101000000000100100100011",
5629 => "0101000110001100101010001",
5630 => "0110000110000100101000011",
5631 => "0010100000001100100110001",
5632 => "0011100000000100100100011",
5633 => "0001000000101010011110001",
5634 => "0100100000001110011100011",
5635 => "0011001011011000010110001",
5636 => "0101001011001000010100011",
5637 => "0100000111010010100010001",
5638 => "0101100111000110100000011",
5639 => "0100100110001101001010001",
5640 => "0100100110000110100100010",
5641 => "0110001111000110100100010",
5642 => "0111101110010000101010001",
5643 => "1001101110001000010100010",
5644 => "0111110011001000010100010",
5645 => "0000101110010000101010001",
5646 => "0000101110001000010100010",
5647 => "0010110011001000010100010",
5648 => "0101100000010000101010001",
5649 => "0111100000001000010100010",
5650 => "0101100101001000010100010",
5651 => "0010100000010000101010001",
5652 => "0010100000001000010100010",
5653 => "0100100101001000010100010",
5654 => "0011000001011000010110001",
5655 => "0011000001001100010100010",
5656 => "0000101100100100001010001",
5657 => "0101001100010010001000010",
5658 => "0001001000101000011010001",
5659 => "0110001000010100001100010",
5660 => "0001001011010100001100010",
5661 => "0011100110010010011110001",
5662 => "0101000110000110011100011",
5663 => "0101000101010001000010001",
5664 => "0111000101001000100000010",
5665 => "0101001101001000100000010",
5666 => "0001101001100000100010001",
5667 => "0001101001010000010000010",
5668 => "0101101101010000010000010",
5669 => "0011101000010100010010001",
5670 => "0011101000001010010000010",
5671 => "0011101100010100100010001",
5672 => "0011101100001010010000010",
5673 => "0110010000001010010000010",
5674 => "0100110011011110010010001",
5675 => "0111010011001010010000011",
5676 => "0000100000100100100110001",
5677 => "0011100000001100100100011",
5678 => "0110100100010100100010001",
5679 => "1001000100001010010000010",
5680 => "0110101000001010010000010",
5681 => "0001110000100100010010001",
5682 => "0100110000001100010000011",
5683 => "0100000111010100110010001",
5684 => "0110100111001010011000010",
5685 => "0100001101001010011000010",
5686 => "0011000111010100110010001",
5687 => "0011000111001010011000010",
5688 => "0101101101001010011000010",
5689 => "0010000110100100011110001",
5690 => "0101000110001100011100011",
5691 => "0000010001100100001110001",
5692 => "0000010010100100000100011",
5693 => "0001110001100100001110001",
5694 => "0001110010100100000100011",
5695 => "0001000100001100101010001",
5696 => "0010000100000100101000011",
5697 => "1000000000010001100010001",
5698 => "1000000000001001100000010",
5699 => "0010000000010000111110001",
5700 => "0100000000001000111100010",
5701 => "1000000000010001100010001",
5702 => "1000000000001001100000010",
5703 => "0000100100100100100110001",
5704 => "0011100100001100100100011",
5705 => "0111101100010010011010001",
5706 => "0111101110010010001000011",
5707 => "0001101001100100011010001",
5708 => "0001101001010010001100010",
5709 => "0110001100010010001100010",
5710 => "1001000101001100100110001",
5711 => "1001001000001100001100011",
5712 => "0000000101001100100110001",
5713 => "0000001000001100001100011",
5714 => "0010000111100100010010001",
5715 => "0110100111010010001000010",
5716 => "0010001001010010001000010",
5717 => "0001000001011001010010001",
5718 => "0001000001001100101000010",
5719 => "0100001011001100101000010",
5720 => "1000100000001101011110001",
5721 => "1000100000000111011100010",
5722 => "0000100110000101001010001",
5723 => "0000101111000100100100010",
5724 => "0100001000010100011010001",
5725 => "0100001010010100001000011",
5726 => "0000000110101000011010001",
5727 => "0000000110010100001100010",
5728 => "0101001001010100001100010",
5729 => "0101101100011000010110001",
5730 => "0111101100001000010100011",
5731 => "0000000100000111001110001",
5732 => "0000100100000011001100011",
5733 => "1001100001000111001010001",
5734 => "1010000001000011001000011",
5735 => "0001000001000111001010001",
5736 => "0001100001000011001000011",
5737 => "0001101010100100001110001",
5738 => "0100101010001100001100011",
5739 => "0010000100010100100110001",
5740 => "0100100100001010100100010",
5741 => "0011101101011100011110001",
5742 => "0011101101001110011100010",
5743 => "0001101101011100011110001",
5744 => "0101001101001110011100010",
5745 => "0100001111010010011010001",
5746 => "0101101111000110011000011",
5747 => "0010001110010000101010001",
5748 => "0010001110001000010100010",
5749 => "0100010011001000010100010",
5750 => "0101001110001000101010001",
5751 => "0101010011001000010100010",
5752 => "0001101000001011000010001",
5753 => "0001110000001010100000010",
5754 => "0111101010010010011010001",
5755 => "0111101100010010001000011",
5756 => "0000001010010010011010001",
5757 => "0000001100010010001000011",
5758 => "0011000111011000100110001",
5759 => "0011001010011000001100011",
5760 => "0100101010001010100010001",
5761 => "0100101110001010010000010",
5762 => "0110000001000110110010001",
5763 => "0110000111000110011000010",
5764 => "0100001111001100100110001",
5765 => "0101001111000100100100011",
5766 => "1000000110001110011010001",
5767 => "1000001001001110001100010",
5768 => "0100000001001001011010001",
5769 => "0101000001000101011000010",
5770 => "0011000110011100001110001",
5771 => "0011000110001110001100010",
5772 => "0000010010100110001110001",
5773 => "0000010011100110000100011",
5774 => "1000100000001101100010001",
5775 => "1000100000000111100000010",
5776 => "0000001101011110011010001",
5777 => "0010101101001010011000011",
5778 => "0100100110010100111010001",
5779 => "0111000110001010011100010",
5780 => "0100101101001010011100010",
5781 => "0000100110010000101010001",
5782 => "0000100110001000010100010",
5783 => "0010101011001000010100010",
5784 => "0011100110011000010110001",
5785 => "0011100110001100010100010",
5786 => "0011100111010010011010001",
5787 => "0101000111000110011000011",
5788 => "0011101000011100111010001",
5789 => "0111001000001110011100010",
5790 => "0011101111001110011100010",
5791 => "0001101000011100111010001",
5792 => "0001101000001110011100010",
5793 => "0101001111001110011100010",
5794 => "0100101000011010010010001",
5795 => "0100101010011010001000010",
5796 => "0001100010001100110010001",
5797 => "0001100010000110011000010",
5798 => "0011001000000110011000010",
5799 => "0011001010100010011010001",
5800 => "0011001101100010001100010",
5801 => "0000101010100010011010001",
5802 => "0000101101100010001100010",
5803 => "1000000111010000100110001",
5804 => "1000001010010000001100011",
5805 => "0000000111010000100110001",
5806 => "0000001010010000001100011",
5807 => "0000001001110000101010001",
5808 => "0110001001011000010100010",
5809 => "0000001110011000010100010",
5810 => "0001100010011110100010001",
5811 => "0100000010001010100000011",
5812 => "0010000010100100100010001",
5813 => "0101000010001100100000011",
5814 => "0000000001100100010010001",
5815 => "0000000001010010001000010",
5816 => "0100100011010010001000010",
5817 => "1010000010000111001010001",
5818 => "1010100010000011001000011",
5819 => "0000100011000111001110001",
5820 => "0001000011000011001100011",
5821 => "1001001000001101000010001",
5822 => "1010001000000101000000011",
5823 => "0000001000001101000010001",
5824 => "0001001000000101000000011",
5825 => "0100010010010110011010001",
5826 => "0100010100010110001000011",
5827 => "0010000110011000010110001",
5828 => "0100000110001000010100011",
5829 => "0011100110011000010110001",
5830 => "0101100110001000010100011",
5831 => "0011000011010010011010001",
5832 => "0100100011000110011000011",
5833 => "0011100110011000010110001",
5834 => "0011100110001100010100010",
5835 => "0100101000001100011110001",
5836 => "0110001000000110011100010",
5837 => "0100000010010010011010001",
5838 => "0101100010000110011000011",
5839 => "0100001110001100100110001",
5840 => "0100010001001100001100011",
5841 => "0100000010010010011010001",
5842 => "0101100010000110011000011",
5843 => "0010000011100001010010001",
5844 => "0010000011010000101000010",
5845 => "0110001101010000101000010",
5846 => "0011100110010100110010001",
5847 => "0110000110001010011000010",
5848 => "0011101100001010011000010",
5849 => "0000000010001110110010001",
5850 => "0000000110001110010000011",
5851 => "0110010001010110011010001",
5852 => "0110010011010110001000011",
5853 => "0010000111011000100010001",
5854 => "0010000111001100010000010",
5855 => "0101001011001100010000010",
5856 => "0100001011010000101010001",
5857 => "0110001011001000010100010",
5858 => "0100010000001000010100010",
5859 => "0100100001001000100110001",
5860 => "0101100001000100100100010",
5861 => "0111000000000111011010001",
5862 => "0111100000000011011000011",
5863 => "0011100000000111011010001",
5864 => "0100000000000011011000011",
5865 => "0010000111100100010010001",
5866 => "0110100111010010001000010",
5867 => "0010001001010010001000010",
5868 => "0101000010001000111110001",
5869 => "0101000111001000010100011",
5870 => "0110000001000110110010001",
5871 => "0110000111000110011000010",
5872 => "0000000000100100110110001",
5873 => "0100100000010010110100010",
5874 => "1000000000000111100010001",
5875 => "1000100000000011100000011",
5876 => "0010100000000111100010001",
5877 => "0011000000000011100000011",
5878 => "0101001111001010100010001",
5879 => "0101010011001010010000010",
5880 => "0001010010100100001010001",
5881 => "0001010011100100000100010",
5882 => "0001001000101000001110001",
5883 => "0001001001101000000100011",
5884 => "0011100110010010011010001",
5885 => "0011101000010010001000011",
5886 => "0001100010100110101010001",
5887 => "0001100111100110010100010",
5888 => "0001000111100110001110001",
5889 => "0001001000100110000100011",
5890 => "0111100110010010010010001",
5891 => "0111101000010010001000010",
5892 => "0001000010100100100010001",
5893 => "0100000010001100100000011",
5894 => "0101001001011100010010001",
5895 => "0101001001001110010000010",
5896 => "0010000100001101000010001",
5897 => "0011100100000111000000010",
5898 => "0111101000010011000010001",
5899 => "1001001000000111000000011",
5900 => "0000001000010011000010001",
5901 => "0001101000000111000000011",
5902 => "1001000000001100111010001",
5903 => "1010000000000100111000011",
5904 => "0000000000001100111010001",
5905 => "0001000000000100111000011",
5906 => "0111100000001101011010001",
5907 => "1000100000000101011000011",
5908 => "0001100000001101011010001",
5909 => "0010100000000101011000011",
5910 => "0110000010011001010010001",
5911 => "1000000010001001010000011",
5912 => "0000000010011001010010001",
5913 => "0010000010001001010000011",
5914 => "0101100110001000100110001",
5915 => "0101100110000100100100010",
5916 => "0100100000001101000010001",
5917 => "0110000000000111000000010",
5918 => "0110000001000110110010001",
5919 => "0110000111000110011000010",
5920 => "0001100100100100011010001",
5921 => "0001100100010010001100010",
5922 => "0110000111010010001100010",
5923 => "0010100101100000100010001",
5924 => "0110100101010000010000010",
5925 => "0010101001010000010000010",
5926 => "0000001101010100011010001",
5927 => "0000001111010100001000011",
5928 => "0100001110010010011010001",
5929 => "0100010000010010001000011",
5930 => "0011000010010010011010001",
5931 => "0100100010000110011000011",
5932 => "0111000001010100100010001",
5933 => "1001100001001010010000010",
5934 => "0111000101001010010000010",
5935 => "0100100001000110110010001",
5936 => "0100100111000110011000010",
5937 => "0011000100011000100110001",
5938 => "0011000111011000001100011",
5939 => "0011000101011000011010001",
5940 => "0101000101001000011000011",
5941 => "0000100001010000010110001",
5942 => "0010100001001000010100010",
5943 => "0110001100001100100010001",
5944 => "0110010000001100010000010",
5945 => "0001101100011000011010001",
5946 => "0001101110011000001000011",
5947 => "0100110010011000011010001",
5948 => "0111110010001100001100010",
5949 => "0100110101001100001100010",
5950 => "0010001101001100011010001",
5951 => "0010010000001100001100010",
5952 => "0101100011001111001010001",
5953 => "0101101100001110100100010",
5954 => "0001101001100100001110001",
5955 => "0100101001001100001100011",
5956 => "0010100011100110001010001",
5957 => "0010100100100110000100010",
5958 => "0010000010011000011010001",
5959 => "0010000010001100001100010",
5960 => "0101000101001100001100010",
5961 => "0100100110001100100110001",
5962 => "0101100110000100100100011",
5963 => "0100000110001100100110001",
5964 => "0101000110000100100100011",
5965 => "1000001001001010111110001",
5966 => "1000001110001010010100011",
5967 => "0001101001001010111110001",
5968 => "0001101110001010010100011",
5969 => "0011000110011100011010001",
5970 => "0110100110001110001100010",
5971 => "0011001001001110001100010",
5972 => "0100000110000110111010001",
5973 => "0100001101000110011100010",
5974 => "0000010000110000010110001",
5975 => "0100010000010000010100011",
5976 => "0000010100101000001110001",
5977 => "0101010100010100001100010",
5978 => "0010101010100100001010001",
5979 => "0010101011100100000100010",
5980 => "0000000110001100101010001",
5981 => "0001000110000100101000011",
5982 => "0001000001101000001110001",
5983 => "0001000010101000000100011",
5984 => "0100101101001100101110001",
5985 => "0101101101000100101100011",
5986 => "0100101111001100100010001",
5987 => "0100110011001100010000010",
5988 => "0100101100001100100110001",
5989 => "0100101111001100001100011",
5990 => "0010101011100100001010001",
5991 => "0010101100100100000100010",
5992 => "0001000110011110011010001",
5993 => "0001001000011110001000011",
5994 => "0011000000100100001110001",
5995 => "0011000001100100000100011",
5996 => "0010100000000111001010001",
5997 => "0011000000000011001000011",
5998 => "1001000011001100101010001",
5999 => "1010000011000100101000011",
6000 => "0000000011001100101010001",
6001 => "0001000011000100101000011",
6002 => "0101000101010000100110001",
6003 => "0101000101001000100100010",
6004 => "0011000101010000100110001",
6005 => "0101000101001000100100010",
6006 => "0001100010101000001110001",
6007 => "0001100011101000000100011",
6008 => "0010100010011010010010001",
6009 => "0010100100011010001000010",
6010 => "1000100000001110111010001",
6011 => "1000100111001110011100010",
6012 => "0000000000001110111010001",
6013 => "0000000111001110011100010",
6014 => "0100101011010100011010001",
6015 => "0100101011001010011000010",
6016 => "0010101011010100011010001",
6017 => "0101001011001010011000010",
6018 => "0101100110000111001010001",
6019 => "0101101100000110011000011",
6020 => "0000010000100100001110001",
6021 => "0000010001100100000100011",
6022 => "0011010000100100001110001",
6023 => "0011010001100100000100011",
6024 => "0010000110010010101010001",
6025 => "0010001011010010010100010",
6026 => "0100100111011110010010001",
6027 => "0100101001011110001000010",
6028 => "0010100110011000011010001",
6029 => "0010100110001100001100010",
6030 => "0101101001001100001100010",
6031 => "0011000001011000100110001",
6032 => "0011000100011000001100011",
6033 => "0011101001001100110010001",
6034 => "0011101001000110011000010",
6035 => "0101001111000110011000010",
6036 => "0101100101011010011010001",
6037 => "0101100111011010001000011",
6038 => "0000101011101100110110001",
6039 => "0110001011010110110100010",
6040 => "1001001000001100011010001",
6041 => "1001001011001100001100010",
6042 => "0000001000001100011010001",
6043 => "0000001011001100001100010",
6044 => "0000000110110000001110001",
6045 => "0000000111110000000100011",
6046 => "0000000101010100011010001",
6047 => "0000000111010100001000011",
6048 => "0011000111100100001110001",
6049 => "0011001000100100000100011",
6050 => "0000000000010100011010001",
6051 => "0000000010010100001000011",
6052 => "1001100000000111001110001",
6053 => "1010000000000011001100011",
6054 => "0010000110011001000010001",
6055 => "0010000110001100100000010",
6056 => "0101001110001100100000010",
6057 => "1001100110001001001010001",
6058 => "1010100110000100100100010",
6059 => "1001101111000100100100010",
6060 => "0000100110001001001010001",
6061 => "0000100110000100100100010",
6062 => "0001101111000100100100010",
6063 => "0001110101100100001110001",
6064 => "0001110110100100000100011",
6065 => "0000010011010010010010001",
6066 => "0000010101010010001000010",
6067 => "0110010010011000011010001",
6068 => "1001010010001100001100010",
6069 => "0110010101001100001100010",
6070 => "0011110010010010010010001",
6071 => "0011110100010010001000010",
6072 => "0110010000010100100010001",
6073 => "1000110000001010010000010",
6074 => "0110010100001010010000010",
6075 => "0001010000010100100010001",
6076 => "0001010000001010010000010",
6077 => "0011110100001010010000010",
6078 => "0111000000010100110010001",
6079 => "1001100000001010011000010",
6080 => "0111000110001010011000010",
6081 => "0000000000010100110010001",
6082 => "0000000000001010011000010",
6083 => "0010100110001010011000010",
6084 => "0111101110010010011010001",
6085 => "0111110000010010001000011",
6086 => "0000001110010010011010001",
6087 => "0000010000010010001000011",
6088 => "0111001110010100011010001",
6089 => "0111010000010100001000011",
6090 => "0000001110010100011010001",
6091 => "0000010000010100001000011",
6092 => "0010110010100100001010001",
6093 => "0010110011100100000100010",
6094 => "0000010010100100001110001",
6095 => "0000010011100100000100011",
6096 => "0001100101100100110010001",
6097 => "0110000101010010011000010",
6098 => "0001101011010010011000010",
6099 => "0010100011001110100110001",
6100 => "0010100110001110001100011",
6101 => "0010000000100110111110001",
6102 => "0010000101100110010100011",
6103 => "0001100000100000010010001",
6104 => "0001100010100000001000010",
6105 => "0010001100100000110010001",
6106 => "0010001100010000110000010",
6107 => "0010000011011000111110001",
6108 => "0101000011001100111100010",
6109 => "1000000100000101001110001",
6110 => "1000000100000011001100010",
6111 => "0011000100000101001110001",
6112 => "0011100100000011001100010",
6113 => "0110101110010000101010001",
6114 => "1000101110001000010100010",
6115 => "0110110011001000010100010",
6116 => "0001101110010000101010001",
6117 => "0001101110001000010100010",
6118 => "0011110011001000010100010",
6119 => "0110000110000111001010001",
6120 => "0110001100000110011000011",
6121 => "0010101011011000011010001",
6122 => "0010101011001100001100010",
6123 => "0101101110001100001100010",
6124 => "0101000101010000101010001",
6125 => "0111000101001000010100010",
6126 => "0101001010001000010100010",
6127 => "0011000100011000101010001",
6128 => "0011000100001100010100010",
6129 => "0110001001001100010100010",
6130 => "0011001000100100101010001",
6131 => "0111101000010010010100010",
6132 => "0011001101010010010100010",
6133 => "0000001000100100101010001",
6134 => "0000001000010010010100010",
6135 => "0100101101010010010100010",
6136 => "0110000110000111001010001",
6137 => "0110001100000110011000011",
6138 => "0000001110100100001110001",
6139 => "0000001111100100000100011",
6140 => "0110000110000111001010001",
6141 => "0110001100000110011000011",
6142 => "0100100110000111001010001",
6143 => "0100101100000110011000011",
6144 => "0011001110100100001110001",
6145 => "0011001111100100000100011",
6146 => "0000000101100100001110001",
6147 => "0000000110100100000100011",
6148 => "0001000101101100001110001",
6149 => "0001000110101100000100011",
6150 => "0000000000101010101010001",
6151 => "0011100000001110101000011",
6152 => "0011000011100101000110001",
6153 => "0110000011001101000100011",
6154 => "0000000011100101000110001",
6155 => "0011000011001101000100011",
6156 => "0000001100110000101110001",
6157 => "0100001100010000101100011",
6158 => "0010001010100000011010001",
6159 => "0010001101100000001100010",
6160 => "0110001000001100100010001",
6161 => "0110001100001100010000010",
6162 => "0011001110010000011110001",
6163 => "0101001110001000011100010",
6164 => "0111101010001100111010001",
6165 => "1001001010000110011100010",
6166 => "0111110001000110011100010",
6167 => "0001101010001100111010001",
6168 => "0001101010000110011100010",
6169 => "0011010001000110011100010",
6170 => "0011001100100100001010001",
6171 => "0011001101100100000100010",
6172 => "0010101000010100011010001",
6173 => "0010101010010100001000011",
6174 => "0110001011010010010010001",
6175 => "0110001101010010001000010",
6176 => "0000001011010010011010001",
6177 => "0000001101010010001000011",
6178 => "0101100010000111001010001",
6179 => "0110000010000011001000011",
6180 => "0101000010000111001010001",
6181 => "0101100010000011001000011",
6182 => "0100101100001100101010001",
6183 => "0101101100000100101000011",
6184 => "0000101010001100100110001",
6185 => "0000101101001100001100011",
6186 => "0011001001100000011010001",
6187 => "0111001001010000001100010",
6188 => "0011001100010000001100010",
6189 => "0000101000010010011010001",
6190 => "0000101010010010001000011",
6191 => "0011100111100000011010001",
6192 => "0011101001100000001000011",
6193 => "0000000000100100001110001",
6194 => "0000000001100100000100011",
6195 => "0101000000001100100110001",
6196 => "0110000000000100100100011",
6197 => "0100100101001100011010001",
6198 => "0110000101000110011000010",
6199 => "0101000110001001001010001",
6200 => "0110000110000100100100010",
6201 => "0101001111000100100100010",
6202 => "0100000000001100100110001",
6203 => "0101000000000100100100011",
6204 => "0100100001001100100110001",
6205 => "0100100100001100001100011",
6206 => "0000100000100100100110001",
6207 => "0000100011100100001100011",
6208 => "0000000011110000001110001",
6209 => "0000000100110000000100011",
6210 => "0011001110010010010010001",
6211 => "0011010000010010001000010",
6212 => "0100001001010000101010001",
6213 => "0110001001001000010100010",
6214 => "0100001110001000010100010",
6215 => "0010100010011010100110001",
6216 => "0010100101011010001100011",
6217 => "0010000100100000100110001",
6218 => "0010000111100000001100011",
6219 => "0010000100011100100110001",
6220 => "0010000111011100001100011",
6221 => "0100000101010010011010001",
6222 => "0100000111010010001000011",
6223 => "0000100111100000011010001",
6224 => "0000101001100000001000011",
6225 => "0101000101011010100110001",
6226 => "0101001000011010001100011",
6227 => "0000100101011010100110001",
6228 => "0000101000011010001100011",
6229 => "0000000100110000011010001",
6230 => "0110000100011000001100010",
6231 => "0000000111011000001100010",
6232 => "0000101110010100100110001",
6233 => "0000110001010100001100011",
6234 => "0010110001100100001110001",
6235 => "0010110010100100000100011",
6236 => "0000010000100100001110001",
6237 => "0000010001100100000100011",
6238 => "0100110001010010011010001",
6239 => "0100110011010010001000011",
6240 => "0000110100101100010010001",
6241 => "0000110100010110001000010",
6242 => "0110010110010110001000010",
6243 => "0100001110010000011010001",
6244 => "0100010001010000001100010",
6245 => "0100000110010000111110001",
6246 => "0100001011010000010100011",
6247 => "0010100100100100001110001",
6248 => "0010100101100100000100011",
6249 => "0100100011001010101010001",
6250 => "0100101000001010010100010",
6251 => "0011001000011000001110001",
6252 => "0011001000001100001100010",
6253 => "0001000110100100011010001",
6254 => "0001000110010010001100010",
6255 => "0101101001010010001100010",
6256 => "0101000110001001001010001",
6257 => "0110000110000100100100010",
6258 => "0101001111000100100100010",
6259 => "0011100101001100011010001",
6260 => "0101000101000110011000010",
6261 => "0111000101000101001010001",
6262 => "0111001110000100100100010",
6263 => "0100000101000101001010001",
6264 => "0100001110000100100100010",
6265 => "0100100010010100011010001",
6266 => "0100100010001010011000010",
6267 => "0001100001100100110010001",
6268 => "0110000001010010110000010",
6269 => "0010100010100011011010001",
6270 => "0010101101100010101100010",
6271 => "0010000000011000011010001",
6272 => "0010000010011000001000011",
6273 => "0011001001100000011010001",
6274 => "0111001001010000001100010",
6275 => "0011001100010000001100010",
6276 => "0100100000001011001010001",
6277 => "0100101001001010100100010",
6278 => "0110000000001100100110001",
6279 => "0111000000000100100100011",
6280 => "0011000000001100100110001",
6281 => "0100000000000100100100011",
6282 => "0100100001001100110010001",
6283 => "0101100001000100110000011",
6284 => "0010101001011010010010001",
6285 => "0010101011011010001000010",
6286 => "0010101000100110001110001",
6287 => "0010101001100110000100011",
6288 => "0100101001001100100010001",
6289 => "0100101101001100010000010",
6290 => "0101101001001000111110001",
6291 => "0101101110001000010100011",
6292 => "0001000000001100111010001",
6293 => "0001000000000110011100010",
6294 => "0010100111000110011100010",
6295 => "0111100001001100111010001",
6296 => "1001000001000110011100010",
6297 => "0111101000000110011100010",
6298 => "0001100001001100111010001",
6299 => "0001100001000110011100010",
6300 => "0011001000000110011100010",
6301 => "0001110100100100010010001",
6302 => "0110010100010010001000010",
6303 => "0001110110010010001000010",
6304 => "0010100000001001010010001",
6305 => "0010100000000100101000010",
6306 => "0011101010000100101000010",
6307 => "1000001000010000110010001",
6308 => "1010001000001000011000010",
6309 => "1000001110001000011000010",
6310 => "0000001000010000110010001",
6311 => "0000001000001000011000010",
6312 => "0010001110001000011000010",
6313 => "0110101101010100100010001",
6314 => "1001001101001010010000010",
6315 => "0110110001001010010000010",
6316 => "0000101101010100100010001",
6317 => "0000101101001010010000010",
6318 => "0011010001001010010000010",
6319 => "0111101000001000111110001",
6320 => "0111101101001000010100011",
6321 => "0010101000001000111110001",
6322 => "0010101101001000010100011",
6323 => "0011001011100000110010001",
6324 => "0011001111100000010000011",
6325 => "0001001011100000110010001",
6326 => "0001001111100000010000011",
6327 => "0111001100001110100110001",
6328 => "0111001111001110001100011",
6329 => "0101000001000111010110001",
6330 => "0101001000000110011100011",
6331 => "0110101011010010010010001",
6332 => "0110101101010010001000010",
6333 => "0001101010100010100110001",
6334 => "0001101101100010001100011",
6335 => "0110101000010000111110001",
6336 => "0110101101010000010100011",
6337 => "0001101000010000111110001",
6338 => "0001101101010000010100011",
6339 => "0101101110010100100010001",
6340 => "1000001110001010010000010",
6341 => "0101110010001010010000010",
6342 => "0000010010101100011010001",
6343 => "0000010010010110001100010",
6344 => "0101110101010110001100010",
6345 => "0000010000110000010010001",
6346 => "0000010000011000010000010",
6347 => "0011010100011000001110001",
6348 => "0110010100001100001100010",
6349 => "1001001100001100110010001",
6350 => "1010101100000110011000010",
6351 => "1001010010000110011000010",
6352 => "0000001100001100110010001",
6353 => "0000001100000110011000010",
6354 => "0001110010000110011000010",
6355 => "0111110001010010011010001",
6356 => "0111110011010010001000011",
6357 => "0000100110101100101010001",
6358 => "0000100110010110010100010",
6359 => "0110001011010110010100010",
6360 => "0111110001010010011010001",
6361 => "0111110011010010001000011",
6362 => "0000010010100100001010001",
6363 => "0000010011100100000100010",
6364 => "0001101111100110001110001",
6365 => "0001110000100110000100011",
6366 => "0000001101100100001110001",
6367 => "0000001110100100000100011",
6368 => "0111110001010010011010001",
6369 => "0111110011010010001000011",
6370 => "0000010001010010011010001",
6371 => "0000010011010010001000011",
6372 => "0110010001010010011010001",
6373 => "0110010011010010001000011",
6374 => "0001110001010010011010001",
6375 => "0001110011010010001000011",
6376 => "1000000010000111010010001",
6377 => "1000100010000011010000011",
6378 => "0000001101110000100010001",
6379 => "0000010001110000010000010",
6380 => "0100100001001101011010001",
6381 => "0110000001000110101100010",
6382 => "0100101100000110101100010"
);

begin

--process for read and write operation.
PROCESS(clk)
BEGIN
    if(rising_edge(clk)) then
        data_o <= ram(adress);
    end if;
END PROCESS;

end Behavioral;

